`timescale 1 ns / 1 ps

module dct_coeff_huffman_decoder (
    input clk,
    input reset,
    input codetable,
    input data_valid,
    input data,
    output bit result_valid,
    output bit [15:0] result
);

    bit [6:0] state;

    typedef struct {
        bit [6:0]  index;  // 0 - 111
        bit [15:0] value;
    } plm_vlc_uint_t;

    // got this from https://github.com/phoboslab/pl_mpeg/blob/master/pl_mpeg.h
    // verilog_format: off

    plm_vlc_uint_t PLM_VIDEO_MACROBLOCK_ADDRESS_INCREMENT[40*2] = '{
        '{  1,    0}, '{  0,    1},  //   0: x
        '{  2,    0}, '{  3,    0},  //   1: 0x
        '{  4,    0}, '{  5,    0},  //   2: 00x
        '{  0,    3}, '{  0,    2},  //   3: 01x
        '{  6,    0}, '{  7,    0},  //   4: 000x
        '{  0,    5}, '{  0,    4},  //   5: 001x
        '{  8,    0}, '{  9,    0},  //   6: 0000x
        '{  0,    7}, '{  0,    6},  //   7: 0001x
        '{ 10,    0}, '{ 11,    0},  //   8: 0000 0x
        '{ 12,    0}, '{ 13,    0},  //   9: 0000 1x
        '{ 14,    0}, '{ 15,    0},  //  10: 0000 00x
        '{ 16,    0}, '{ 17,    0},  //  11: 0000 01x
        '{ 18,    0}, '{ 19,    0},  //  12: 0000 10x
        '{  0,    9}, '{  0,    8},  //  13: 0000 11x
        '{  0,    0}, '{ 20,    0},  //  14: 0000 000x
        '{  0,    0}, '{ 21,    0},  //  15: 0000 001x
        '{ 22,    0}, '{ 23,    0},  //  16: 0000 010x
        '{  0,   15}, '{  0,   14},  //  17: 0000 011x
        '{  0,   13}, '{  0,   12},  //  18: 0000 100x
        '{  0,   11}, '{  0,   10},  //  19: 0000 101x
        '{ 24,    0}, '{ 25,    0},  //  20: 0000 0001x
        '{ 26,    0}, '{ 27,    0},  //  21: 0000 0011x
        '{ 28,    0}, '{ 29,    0},  //  22: 0000 0100x
        '{ 30,    0}, '{ 31,    0},  //  23: 0000 0101x
        '{ 32,    0}, '{  0,    0},  //  24: 0000 0001 0x
        '{  0,    0}, '{ 33,    0},  //  25: 0000 0001 1x
        '{ 34,    0}, '{ 35,    0},  //  26: 0000 0011 0x
        '{ 36,    0}, '{ 37,    0},  //  27: 0000 0011 1x
        '{ 38,    0}, '{ 39,    0},  //  28: 0000 0100 0x
        '{  0,   21}, '{  0,   20},  //  29: 0000 0100 1x
        '{  0,   19}, '{  0,   18},  //  30: 0000 0101 0x
        '{  0,   17}, '{  0,   16},  //  31: 0000 0101 1x
        '{  0,   35}, '{  0,    0},  //  32: 0000 0001 00x
        '{  0,    0}, '{  0,   34},  //  33: 0000 0001 11x
        '{  0,   33}, '{  0,   32},  //  34: 0000 0011 00x
        '{  0,   31}, '{  0,   30},  //  35: 0000 0011 01x
        '{  0,   29}, '{  0,   28},  //  36: 0000 0011 10x
        '{  0,   27}, '{  0,   26},  //  37: 0000 0011 11x
        '{  0,   25}, '{  0,   24},  //  38: 0000 0100 00x
        '{  0,   23}, '{  0,   22}   //  39: 0000 0100 01x
    };

    plm_vlc_uint_t PLM_VIDEO_DCT_COEFF[112*2] = '{
        '{   1,        0}, '{   0, 16'h0001},  //   0: x
        '{   2,        0}, '{   3,        0},  //   1: 0x
        '{   4,        0}, '{   5,        0},  //   2: 00x
        '{   6,        0}, '{   0, 16'h0101},  //   3: 01x
        '{   7,        0}, '{   8,        0},  //   4: 000x
        '{   9,        0}, '{  10,        0},  //   5: 001x
        '{   0, 16'h0002}, '{   0, 16'h0201},  //   6: 010x
        '{  11,        0}, '{  12,        0},  //   7: 0000x
        '{  13,        0}, '{  14,        0},  //   8: 0001x
        '{  15,        0}, '{   0, 16'h0003},  //   9: 0010x
        '{   0, 16'h0401}, '{   0, 16'h0301},  //  10: 0011x
        '{  16,        0}, '{   0, 16'hffff},  //  11: 0000 0x
        '{  17,        0}, '{  18,        0},  //  12: 0000 1x
        '{   0, 16'h0701}, '{   0, 16'h0601},  //  13: 0001 0x
        '{   0, 16'h0102}, '{   0, 16'h0501},  //  14: 0001 1x
        '{  19,        0}, '{  20,        0},  //  15: 0010 0x
        '{  21,        0}, '{  22,        0},  //  16: 0000 00x
        '{   0, 16'h0202}, '{   0, 16'h0901},  //  17: 0000 10xw
        '{   0, 16'h0004}, '{   0, 16'h0801},  //  18: 0000 11x
        '{  23,        0}, '{  24,        0},  //  19: 0010 00x
        '{  25,        0}, '{  26,        0},  //  20: 0010 01x
        '{  27,        0}, '{  28,        0},  //  21: 0000 000x
        '{  29,        0}, '{  30,        0},  //  22: 0000 001x
        '{   0, 16'h0d01}, '{   0, 16'h0006},  //  23: 0010 000x
        '{   0, 16'h0c01}, '{   0, 16'h0b01},  //  24: 0010 001x
        '{   0, 16'h0302}, '{   0, 16'h0103},  //  25: 0010 010x
        '{   0, 16'h0005}, '{   0, 16'h0a01},  //  26: 0010 011x
        '{  31,        0}, '{  32,        0},  //  27: 0000 0000x
        '{  33,        0}, '{  34,        0},  //  28: 0000 0001x
        '{  35,        0}, '{  36,        0},  //  29: 0000 0010x
        '{  37,        0}, '{  38,        0},  //  30: 0000 0011x
        '{  39,        0}, '{  40,        0},  //  31: 0000 0000 0x
        '{  41,        0}, '{  42,        0},  //  32: 0000 0000 1x
        '{  43,        0}, '{  44,        0},  //  33: 0000 0001 0x
        '{  45,        0}, '{  46,        0},  //  34: 0000 0001 1x
        '{   0, 16'h1001}, '{   0, 16'h0502},  //  35: 0000 0010 0x
        '{   0, 16'h0007}, '{   0, 16'h0203},  //  36: 0000 0010 1x
        '{   0, 16'h0104}, '{   0, 16'h0f01},  //  37: 0000 0011 0x
        '{   0, 16'h0e01}, '{   0, 16'h0402},  //  38: 0000 0011 1x
        '{  47,        0}, '{  48,        0},  //  39: 0000 0000 00x
        '{  49,        0}, '{  50,        0},  //  40: 0000 0000 01x
        '{  51,        0}, '{  52,        0},  //  41: 0000 0000 10x
        '{  53,        0}, '{  54,        0},  //  42: 0000 0000 11x
        '{  55,        0}, '{  56,        0},  //  43: 0000 0001 00x
        '{  57,        0}, '{  58,        0},  //  44: 0000 0001 01x
        '{  59,        0}, '{  60,        0},  //  45: 0000 0001 10x
        '{  61,        0}, '{  62,        0},  //  46: 0000 0001 11x
        '{   0,        0}, '{  63,        0},  //  47: 0000 0000 000x
        '{  64,        0}, '{  65,        0},  //  48: 0000 0000 001x
        '{  66,        0}, '{  67,        0},  //  49: 0000 0000 010x
        '{  68,        0}, '{  69,        0},  //  50: 0000 0000 011x
        '{  70,        0}, '{  71,        0},  //  51: 0000 0000 100x
        '{  72,        0}, '{  73,        0},  //  52: 0000 0000 101x
        '{  74,        0}, '{  75,        0},  //  53: 0000 0000 110x
        '{  76,        0}, '{  77,        0},  //  54: 0000 0000 111x
        '{   0, 16'h000b}, '{   0, 16'h0802},  //  55: 0000 0001 000x
        '{   0, 16'h0403}, '{   0, 16'h000a},  //  56: 0000 0001 001x
        '{   0, 16'h0204}, '{   0, 16'h0702},  //  57: 0000 0001 010x
        '{   0, 16'h1501}, '{   0, 16'h1401},  //  58: 0000 0001 011x
        '{   0, 16'h0009}, '{   0, 16'h1301},  //  59: 0000 0001 100x
        '{   0, 16'h1201}, '{   0, 16'h0105},  //  60: 0000 0001 101x
        '{   0, 16'h0303}, '{   0, 16'h0008},  //  61: 0000 0001 110x
        '{   0, 16'h0602}, '{   0, 16'h1101},  //  62: 0000 0001 111x
        '{  78,        0}, '{  79,        0},  //  63: 0000 0000 0001x
        '{  80,        0}, '{  81,        0},  //  64: 0000 0000 0010x
        '{  82,        0}, '{  83,        0},  //  65: 0000 0000 0011x
        '{  84,        0}, '{  85,        0},  //  66: 0000 0000 0100x
        '{  86,        0}, '{  87,        0},  //  67: 0000 0000 0101x
        '{  88,        0}, '{  89,        0},  //  68: 0000 0000 0110x
        '{  90,        0}, '{  91,        0},  //  69: 0000 0000 0111x
        '{   0, 16'h0a02}, '{   0, 16'h0902},  //  70: 0000 0000 1000x
        '{   0, 16'h0503}, '{   0, 16'h0304},  //  71: 0000 0000 1001x
        '{   0, 16'h0205}, '{   0, 16'h0107},  //  72: 0000 0000 1010x
        '{   0, 16'h0106}, '{   0, 16'h000f},  //  73: 0000 0000 1011x
        '{   0, 16'h000e}, '{   0, 16'h000d},  //  74: 0000 0000 1100x
        '{   0, 16'h000c}, '{   0, 16'h1a01},  //  75: 0000 0000 1101x
        '{   0, 16'h1901}, '{   0, 16'h1801},  //  76: 0000 0000 1110x
        '{   0, 16'h1701}, '{   0, 16'h1601},  //  77: 0000 0000 1111x
        '{  92,        0}, '{  93,        0},  //  78: 0000 0000 0001 0x
        '{  94,        0}, '{  95,        0},  //  79: 0000 0000 0001 1x
        '{  96,        0}, '{  97,        0},  //  80: 0000 0000 0010 0x
        '{  98,        0}, '{  99,        0},  //  81: 0000 0000 0010 1x
        '{ 100,        0}, '{ 101,        0},  //  82: 0000 0000 0011 0x
        '{ 102,        0}, '{ 103,        0},  //  83: 0000 0000 0011 1x
        '{   0, 16'h001f}, '{   0, 16'h001e},  //  84: 0000 0000 0100 0x
        '{   0, 16'h001d}, '{   0, 16'h001c},  //  85: 0000 0000 0100 1x
        '{   0, 16'h001b}, '{   0, 16'h001a},  //  86: 0000 0000 0101 0x
        '{   0, 16'h0019}, '{   0, 16'h0018},  //  87: 0000 0000 0101 1x
        '{   0, 16'h0017}, '{   0, 16'h0016},  //  88: 0000 0000 0110 0x
        '{   0, 16'h0015}, '{   0, 16'h0014},  //  89: 0000 0000 0110 1x
        '{   0, 16'h0013}, '{   0, 16'h0012},  //  90: 0000 0000 0111 0x
        '{   0, 16'h0011}, '{   0, 16'h0010},  //  91: 0000 0000 0111 1x
        '{ 104,        0}, '{ 105,        0},  //  92: 0000 0000 0001 00x
        '{ 106,        0}, '{ 107,        0},  //  93: 0000 0000 0001 01x
        '{ 108,        0}, '{ 109,        0},  //  94: 0000 0000 0001 10x
        '{ 110,        0}, '{ 111,        0},  //  95: 0000 0000 0001 11x
        '{   0, 16'h0028}, '{   0, 16'h0027},  //  96: 0000 0000 0010 00x
        '{   0, 16'h0026}, '{   0, 16'h0025},  //  97: 0000 0000 0010 01x
        '{   0, 16'h0024}, '{   0, 16'h0023},  //  98: 0000 0000 0010 10x
        '{   0, 16'h0022}, '{   0, 16'h0021},  //  99: 0000 0000 0010 11x
        '{   0, 16'h0020}, '{   0, 16'h010e},  // 100: 0000 0000 0011 00x
        '{   0, 16'h010d}, '{   0, 16'h010c},  // 101: 0000 0000 0011 01x
        '{   0, 16'h010b}, '{   0, 16'h010a},  // 102: 0000 0000 0011 10x
        '{   0, 16'h0109}, '{   0, 16'h0108},  // 103: 0000 0000 0011 11x
        '{   0, 16'h0112}, '{   0, 16'h0111},  // 104: 0000 0000 0001 000x
        '{   0, 16'h0110}, '{   0, 16'h010f},  // 105: 0000 0000 0001 001x
        '{   0, 16'h0603}, '{   0, 16'h1002},  // 106: 0000 0000 0001 010x
        '{   0, 16'h0f02}, '{   0, 16'h0e02},  // 107: 0000 0000 0001 011x
        '{   0, 16'h0d02}, '{   0, 16'h0c02},  // 108: 0000 0000 0001 100x
        '{   0, 16'h0b02}, '{   0, 16'h1f01},  // 109: 0000 0000 0001 101x
        '{   0, 16'h1e01}, '{   0, 16'h1d01},  // 110: 0000 0000 0001 110x
        '{   0, 16'h1c01}, '{   0, 16'h1b01}   // 111: 0000 0000 0001 111x
    };
    // verilog_format: on

    plm_vlc_uint_t current_entry;
    wire reached_final_state = current_entry.index == 0;

    always_comb begin
        if (codetable) current_entry = PLM_VIDEO_MACROBLOCK_ADDRESS_INCREMENT[{state[5:0], data}];
        else current_entry = PLM_VIDEO_DCT_COEFF[{state, data}];
    end

    always_ff @(posedge clk) begin
        result_valid <= 0;

        if (reset) begin
            state <= 0;
        end else if (data_valid) begin
            if (reached_final_state) begin
                result_valid <= 1;
                result <= current_entry.value;
                state <= 0;
            end else begin
                state <= current_entry.index;
            end
        end
    end

endmodule
