// verilator lint_off UNOPTFLAT
// verilator lint_off INITIALDLY
// verilator lint_off COMBDLY
// verilator lint_off CASEINCOMPLETE
// verilator lint_off UNSIGNED
// verilator lint_off LATCH

module tg68k_alu_2_0_2_0
  (input  clk,
   input  reset,
   input  clkena_lw,
   input  [1:0] cpu,
   input  execopc,
   input  decodeopc,
   input  exe_condition,
   input  exec_tas,
   input  long_start,
   input  non_aligned,
   input  check_aligned,
   input  movem_presub,
   input  set_stop,
   input  z_error,
   input  [1:0] rot_bits,
   input  [88:0] exec,
   input  [31:0] op1out,
   input  [31:0] op2out,
   input  [31:0] reg_qa,
   input  [31:0] reg_qb,
   input  [15:0] opcode,
   input  [15:0] exe_opcode,
   input  [1:0] exe_datatype,
   input  [15:0] sndopc,
   input  [15:0] last_data_read,
   input  [15:0] data_read,
   input  [7:0] flagssr,
   input  [6:0] micro_state,
   input  [7:0] bf_ext_in,
   input  [5:0] bf_shift,
   input  [5:0] bf_width,
   input  [31:0] bf_ffo_offset,
   input  [4:0] bf_loffset,
   output [7:0] bf_ext_out,
   output set_v_flag,
   output [7:0] flags,
   output [2:0] c_out,
   output [31:0] addsub_q,
   output [31:0] aluout);
  wire [31:0] op1in;
  wire [31:0] addsub_a;
  wire [31:0] addsub_b;
  wire [33:0] notaddsub_b;
  wire [33:0] add_result;
  wire [2:0] addsub_ofl;
  wire opaddsub;
  wire [3:0] c_in;
  wire [2:0] flag_z;
  wire [3:0] set_flags;
  wire [7:0] ccrin;
  wire [3:0] last_flags1;
  wire [9:0] bcd_pur;
  wire [8:0] bcd_kor;
  wire halve_carry;
  wire vflag_a;
  wire bcd_a_carry;
  wire [8:0] bcd_a;
  wire [127:0] result_mulu;
  wire [63:0] result_div;
  wire [31:0] result_div_pre;
  wire set_mv_flag;
  wire v_flag;
  wire rot_rot;
  wire rot_lsb;
  wire rot_msb;
  wire rot_x;
  wire rot_c;
  wire [31:0] rot_out;
  wire asl_vflag;
  wire [4:0] bit_number;
  wire [31:0] bits_out;
  wire one_bit_in;
  wire bchg;
  wire bset;
  wire mulu_sign;
  wire muls_msb;
  wire [63:0] mulu_reg;
  wire fasign;
  wire [31:0] faktorb;
  wire [63:0] div_reg;
  wire [63:0] div_quot;
  wire div_neg;
  wire div_bit;
  wire [32:0] div_sub;
  wire [32:0] div_over;
  wire nozero;
  wire div_qsign;
  wire [63:0] dividend;
  wire divs;
  wire signedop;
  wire op1_sign;
  wire [15:0] op2outext;
  wire [31:0] datareg;
  wire [31:0] bf_datareg;
  wire [39:0] result;
  wire [39:0] result_tmp;
  wire [31:0] unshifted_bitmask;
  wire [39:0] inmux0;
  wire [39:0] inmux1;
  wire [39:0] inmux2;
  wire [31:0] inmux3;
  wire [39:0] shifted_bitmask;
  wire [37:0] bitmaskmux0;
  wire [35:0] bitmaskmux1;
  wire [31:0] bitmaskmux2;
  wire [31:0] bitmaskmux3;
  wire [31:0] bf_set2;
  wire [39:0] shift;
  wire [5:0] bf_firstbit;
  wire [3:0] mux;
  wire [4:0] bitnr;
  wire [31:0] mask;
  wire mask_not_zero;
  wire bf_bset;
  wire bf_nflag;
  wire bf_bchg;
  wire bf_ins;
  wire bf_exts;
  wire bf_fffo;
  wire bf_d32;
  wire bf_s32;
  wire [33:0] hot_msb;
  wire [32:0] vector;
  wire [65:0] result_bs;
  wire [5:0] bit_nr;
  wire [5:0] bit_msb;
  wire [5:0] bs_shift;
  wire [5:0] bs_shift_mod;
  wire [32:0] asl_over;
  wire [32:0] asl_over_xor;
  wire [32:0] asr_sign;
  wire msb;
  wire [5:0] ring;
  wire [31:0] alu;
  wire [31:0] bsout;
  wire bs_v;
  wire bs_c;
  wire bs_x;
  wire n9794_o;
  wire n9795_o;
  wire [23:0] n9796_o;
  wire [6:0] n9797_o;
  wire n9798_o;
  wire [31:0] n9799_o;
  wire [31:0] n9800_o;
  wire [31:0] n9801_o;
  wire [31:0] n9802_o;
  wire [31:0] n9803_o;
  wire [31:0] n9804_o;
  wire n9805_o;
  wire n9806_o;
  wire n9807_o;
  wire [7:0] n9808_o;
  wire n9809_o;
  wire n9811_o;
  wire n9812_o;
  wire n9814_o;
  wire [31:0] n9815_o;
  wire [31:0] n9816_o;
  wire [31:0] n9817_o;
  wire n9818_o;
  wire n9820_o;
  wire n9821_o;
  wire n9823_o;
  wire [15:0] n9824_o;
  wire [15:0] n9825_o;
  wire [31:0] n9826_o;
  wire n9827_o;
  wire [31:0] n9828_o;
  wire [31:0] n9829_o;
  wire [31:0] n9830_o;
  wire [31:0] n9831_o;
  wire n9832_o;
  wire [31:0] n9833_o;
  wire n9834_o;
  wire [31:0] n9835_o;
  wire n9836_o;
  wire [3:0] n9837_o;
  wire [3:0] n9838_o;
  wire [7:0] n9839_o;
  wire n9840_o;
  wire [31:0] n9841_o;
  wire n9842_o;
  wire n9843_o;
  wire n9844_o;
  wire n9845_o;
  wire [15:0] n9846_o;
  wire [15:0] n9847_o;
  wire [31:0] n9848_o;
  wire n9849_o;
  wire n9850_o;
  wire n9851_o;
  wire n9852_o;
  wire [7:0] n9854_o;
  wire n9855_o;
  wire [3:0] n9856_o;
  wire [3:0] n9857_o;
  wire [7:0] n9858_o;
  wire [7:0] n9859_o;
  wire [7:0] n9860_o;
  wire [15:0] n9861_o;
  wire [7:0] n9862_o;
  wire [7:0] n9863_o;
  wire [7:0] n9864_o;
  wire [7:0] n9865_o;
  wire [7:0] n9866_o;
  wire [15:0] n9867_o;
  wire [15:0] n9868_o;
  wire [15:0] n9869_o;
  wire [15:0] n9870_o;
  wire [15:0] n9871_o;
  wire [15:0] n9872_o;
  wire [31:0] n9873_o;
  wire [31:0] n9874_o;
  wire [31:0] n9875_o;
  wire [31:0] n9876_o;
  wire [31:0] n9877_o;
  wire [31:0] n9878_o;
  wire [31:0] n9879_o;
  wire [7:0] n9880_o;
  wire [7:0] n9881_o;
  wire [23:0] n9882_o;
  wire [23:0] n9883_o;
  wire [23:0] n9884_o;
  wire [31:0] n9885_o;
  wire [31:0] n9886_o;
  wire [31:0] n9887_o;
  wire [31:0] n9888_o;
  wire [31:0] n9889_o;
  wire [7:0] n9890_o;
  wire [7:0] n9891_o;
  wire [23:0] n9892_o;
  wire [23:0] n9893_o;
  wire [23:0] n9894_o;
  wire n9899_o;
  wire n9900_o;
  wire n9901_o;
  wire n9902_o;
  wire [1:0] n9903_o;
  wire n9904_o;
  wire [2:0] n9905_o;
  wire [28:0] n9906_o;
  wire [31:0] n9907_o;
  wire [1:0] n9908_o;
  wire [31:0] n9910_o;
  wire [31:0] n9911_o;
  wire [31:0] n9912_o;
  wire n9913_o;
  wire n9916_o;
  wire n9918_o;
  wire [3:0] n9919_o;
  wire [7:0] n9921_o;
  wire [11:0] n9923_o;
  wire [3:0] n9924_o;
  wire [15:0] n9925_o;
  wire n9926_o;
  wire n9927_o;
  wire n9928_o;
  wire n9929_o;
  wire n9930_o;
  wire n9931_o;
  wire n9932_o;
  wire n9933_o;
  wire n9935_o;
  wire n9936_o;
  wire n9937_o;
  wire n9938_o;
  wire n9939_o;
  wire n9940_o;
  wire n9942_o;
  wire n9943_o;
  wire n9944_o;
  wire n9945_o;
  wire n9946_o;
  wire n9947_o;
  wire n9948_o;
  wire n9949_o;
  wire [31:0] n9952_o;
  wire [31:0] n9954_o;
  wire [31:0] n9956_o;
  wire n9957_o;
  wire n9958_o;
  wire n9959_o;
  wire n9960_o;
  wire n9961_o;
  wire n9963_o;
  wire n9964_o;
  wire [31:0] n9965_o;
  wire n9966_o;
  wire n9967_o;
  wire [15:0] n9968_o;
  wire [15:0] n9969_o;
  wire [15:0] n9970_o;
  wire [15:0] n9971_o;
  wire [15:0] n9972_o;
  wire n9974_o;
  wire n9975_o;
  wire n9976_o;
  wire n9977_o;
  wire n9978_o;
  wire n9979_o;
  wire n9980_o;
  wire [31:0] n9982_o;
  wire [31:0] n9983_o;
  wire n9984_o;
  wire n9985_o;
  wire n9987_o;
  wire [31:0] n9990_o;
  wire [31:0] n9991_o;
  wire [31:0] n9992_o;
  wire [31:0] n9993_o;
  wire [31:0] n9994_o;
  wire [31:0] n9995_o;
  wire n9996_o;
  wire n9997_o;
  wire [32:0] n9999_o;
  wire n10000_o;
  wire [33:0] n10001_o;
  wire [32:0] n10003_o;
  wire n10004_o;
  wire [33:0] n10005_o;
  wire [33:0] n10006_o;
  wire [33:0] n10007_o;
  wire [32:0] n10009_o;
  wire n10010_o;
  wire [33:0] n10011_o;
  wire [33:0] n10012_o;
  wire n10013_o;
  wire n10014_o;
  wire n10015_o;
  wire n10016_o;
  wire n10017_o;
  wire n10018_o;
  wire n10019_o;
  wire n10020_o;
  wire n10021_o;
  wire n10022_o;
  wire n10023_o;
  wire [31:0] n10024_o;
  wire n10025_o;
  wire n10026_o;
  wire n10027_o;
  wire n10028_o;
  wire n10029_o;
  wire n10030_o;
  wire n10031_o;
  wire n10032_o;
  wire n10033_o;
  wire n10034_o;
  wire n10035_o;
  wire n10036_o;
  wire n10037_o;
  wire n10038_o;
  wire n10039_o;
  wire n10040_o;
  wire n10041_o;
  wire n10042_o;
  wire n10043_o;
  wire n10044_o;
  wire n10045_o;
  wire [2:0] n10046_o;
  wire n10050_o;
  wire [8:0] n10051_o;
  wire [9:0] n10052_o;
  wire n10053_o;
  wire n10054_o;
  wire n10055_o;
  wire n10056_o;
  wire n10057_o;
  wire [3:0] n10060_o;
  localparam [8:0] n10061_o = 9'b000000000;
  wire n10063_o;
  wire [3:0] n10065_o;
  wire [3:0] n10066_o;
  wire n10067_o;
  wire n10068_o;
  wire n10069_o;
  wire n10070_o;
  wire n10071_o;
  wire n10072_o;
  wire [8:0] n10073_o;
  wire [8:0] n10074_o;
  wire n10075_o;
  wire n10076_o;
  wire n10077_o;
  wire n10078_o;
  wire n10079_o;
  wire [3:0] n10081_o;
  wire n10082_o;
  wire n10083_o;
  wire n10084_o;
  wire n10085_o;
  wire n10086_o;
  wire n10087_o;
  wire n10088_o;
  wire n10089_o;
  wire n10090_o;
  wire n10091_o;
  wire n10092_o;
  wire n10093_o;
  wire n10094_o;
  wire [3:0] n10096_o;
  wire n10097_o;
  wire n10098_o;
  wire n10099_o;
  wire n10100_o;
  wire [8:0] n10101_o;
  wire [8:0] n10102_o;
  wire [7:0] n10103_o;
  wire [7:0] n10104_o;
  wire [7:0] n10105_o;
  wire n10106_o;
  wire [8:0] n10107_o;
  wire n10108_o;
  wire n10110_o;
  wire n10111_o;
  wire n10112_o;
  wire n10113_o;
  wire [1:0] n10118_o;
  wire n10120_o;
  wire n10122_o;
  wire [1:0] n10123_o;
  reg n10126_o;
  reg n10130_o;
  wire n10136_o;
  wire n10137_o;
  wire [1:0] n10138_o;
  wire n10140_o;
  wire [4:0] n10141_o;
  wire [2:0] n10142_o;
  wire [4:0] n10144_o;
  wire [4:0] n10145_o;
  wire [1:0] n10146_o;
  wire n10148_o;
  wire [4:0] n10149_o;
  wire [2:0] n10150_o;
  wire [4:0] n10152_o;
  wire [4:0] n10153_o;
  wire [4:0] n10154_o;
  wire n10160_o;
  wire n10161_o;
  wire n10162_o;
  wire [1:0] n10168_o;
  wire n10170_o;
  wire n10173_o;
  wire [2:0] n10175_o;
  wire n10177_o;
  wire n10179_o;
  wire n10181_o;
  wire n10183_o;
  wire n10185_o;
  wire [4:0] n10186_o;
  reg n10189_o;
  reg n10193_o;
  reg n10197_o;
  reg n10201_o;
  reg n10205_o;
  reg n10208_o;
  wire [1:0] n10209_o;
  wire n10211_o;
  wire n10214_o;
  wire [7:0] n10216_o;
  wire [4:0] n10234_o;
  wire n10236_o;
  wire n10239_o;
  wire n10240_o;
  wire n10241_o;
  wire n10242_o;
  wire n10247_o;
  localparam [31:0] n10248_o = 32'b00000000000000000000000000000000;
  wire [4:0] n10250_o;
  wire n10252_o;
  wire n10255_o;
  wire n10256_o;
  wire n10257_o;
  wire n10258_o;
  wire n10262_o;
  wire n10263_o;
  wire [4:0] n10265_o;
  wire n10267_o;
  wire n10270_o;
  wire n10271_o;
  wire n10272_o;
  wire n10273_o;
  wire n10277_o;
  wire n10278_o;
  wire [4:0] n10280_o;
  wire n10282_o;
  wire n10285_o;
  wire n10286_o;
  wire n10287_o;
  wire n10288_o;
  wire n10292_o;
  wire n10293_o;
  wire [4:0] n10295_o;
  wire n10297_o;
  wire n10300_o;
  wire n10301_o;
  wire n10302_o;
  wire n10303_o;
  wire n10307_o;
  wire n10308_o;
  wire [4:0] n10310_o;
  wire n10312_o;
  wire n10315_o;
  wire n10316_o;
  wire n10317_o;
  wire n10318_o;
  wire n10322_o;
  wire n10323_o;
  wire [4:0] n10325_o;
  wire n10327_o;
  wire n10330_o;
  wire n10331_o;
  wire n10332_o;
  wire n10333_o;
  wire n10337_o;
  wire n10338_o;
  wire [4:0] n10340_o;
  wire n10342_o;
  wire n10345_o;
  wire n10346_o;
  wire n10347_o;
  wire n10348_o;
  wire n10352_o;
  wire n10353_o;
  wire [4:0] n10355_o;
  wire n10357_o;
  wire n10360_o;
  wire n10361_o;
  wire n10362_o;
  wire n10363_o;
  wire n10367_o;
  wire n10368_o;
  wire [4:0] n10370_o;
  wire n10372_o;
  wire n10375_o;
  wire n10376_o;
  wire n10377_o;
  wire n10378_o;
  wire n10382_o;
  wire n10383_o;
  wire [4:0] n10385_o;
  wire n10387_o;
  wire n10390_o;
  wire n10391_o;
  wire n10392_o;
  wire n10393_o;
  wire n10397_o;
  wire n10398_o;
  wire [4:0] n10400_o;
  wire n10402_o;
  wire n10405_o;
  wire n10406_o;
  wire n10407_o;
  wire n10408_o;
  wire n10412_o;
  wire n10413_o;
  wire [4:0] n10415_o;
  wire n10417_o;
  wire n10420_o;
  wire n10421_o;
  wire n10422_o;
  wire n10423_o;
  wire n10427_o;
  wire n10428_o;
  wire [4:0] n10430_o;
  wire n10432_o;
  wire n10435_o;
  wire n10436_o;
  wire n10437_o;
  wire n10438_o;
  wire n10442_o;
  wire n10443_o;
  wire [4:0] n10445_o;
  wire n10447_o;
  wire n10450_o;
  wire n10451_o;
  wire n10452_o;
  wire n10453_o;
  wire n10457_o;
  wire n10458_o;
  wire [4:0] n10460_o;
  wire n10462_o;
  wire n10465_o;
  wire n10466_o;
  wire n10467_o;
  wire n10468_o;
  wire n10472_o;
  wire n10473_o;
  wire [4:0] n10475_o;
  wire n10477_o;
  wire n10480_o;
  wire n10481_o;
  wire n10482_o;
  wire n10483_o;
  wire n10487_o;
  wire n10488_o;
  wire [4:0] n10490_o;
  wire n10492_o;
  wire n10495_o;
  wire n10496_o;
  wire n10497_o;
  wire n10498_o;
  wire n10502_o;
  wire n10503_o;
  wire [4:0] n10505_o;
  wire n10507_o;
  wire n10510_o;
  wire n10511_o;
  wire n10512_o;
  wire n10513_o;
  wire n10517_o;
  wire n10518_o;
  wire [4:0] n10520_o;
  wire n10522_o;
  wire n10525_o;
  wire n10526_o;
  wire n10527_o;
  wire n10528_o;
  wire n10532_o;
  wire n10533_o;
  wire [4:0] n10535_o;
  wire n10537_o;
  wire n10540_o;
  wire n10541_o;
  wire n10542_o;
  wire n10543_o;
  wire n10547_o;
  wire n10548_o;
  wire [4:0] n10550_o;
  wire n10552_o;
  wire n10555_o;
  wire n10556_o;
  wire n10557_o;
  wire n10558_o;
  wire n10562_o;
  wire n10563_o;
  wire [4:0] n10565_o;
  wire n10567_o;
  wire n10570_o;
  wire n10571_o;
  wire n10572_o;
  wire n10573_o;
  wire n10577_o;
  wire n10578_o;
  wire [4:0] n10580_o;
  wire n10582_o;
  wire n10585_o;
  wire n10586_o;
  wire n10587_o;
  wire n10588_o;
  wire n10592_o;
  wire n10593_o;
  wire [4:0] n10595_o;
  wire n10597_o;
  wire n10600_o;
  wire n10601_o;
  wire n10602_o;
  wire n10603_o;
  wire n10607_o;
  wire n10608_o;
  wire [4:0] n10610_o;
  wire n10612_o;
  wire n10615_o;
  wire n10616_o;
  wire n10617_o;
  wire n10618_o;
  wire n10622_o;
  wire n10623_o;
  wire [4:0] n10625_o;
  wire n10627_o;
  wire n10630_o;
  wire n10631_o;
  wire n10632_o;
  wire n10633_o;
  wire n10637_o;
  wire n10638_o;
  wire [4:0] n10640_o;
  wire n10642_o;
  wire n10645_o;
  wire n10646_o;
  wire n10647_o;
  wire n10648_o;
  wire n10652_o;
  wire n10653_o;
  wire [4:0] n10655_o;
  wire n10657_o;
  wire n10660_o;
  wire n10661_o;
  wire n10662_o;
  wire n10663_o;
  wire n10667_o;
  wire n10668_o;
  wire [4:0] n10670_o;
  wire n10672_o;
  wire n10675_o;
  wire n10676_o;
  wire n10677_o;
  wire n10678_o;
  wire n10682_o;
  wire n10683_o;
  wire [4:0] n10685_o;
  wire n10687_o;
  wire n10690_o;
  wire n10691_o;
  wire n10692_o;
  wire n10693_o;
  wire n10694_o;
  wire n10695_o;
  wire n10696_o;
  wire n10697_o;
  wire n10698_o;
  wire n10699_o;
  wire [4:0] n10700_o;
  wire n10702_o;
  wire n10705_o;
  wire n10706_o;
  wire [4:0] n10708_o;
  wire n10711_o;
  wire [31:0] n10712_o;
  wire [31:0] n10713_o;
  wire n10714_o;
  wire [15:0] n10715_o;
  wire [15:0] n10716_o;
  wire [31:0] n10717_o;
  wire [31:0] n10718_o;
  wire n10719_o;
  wire [23:0] n10720_o;
  wire [7:0] n10721_o;
  wire [31:0] n10722_o;
  wire [31:0] n10723_o;
  wire n10724_o;
  wire [35:0] n10726_o;
  wire [3:0] n10727_o;
  wire [3:0] n10728_o;
  wire [3:0] n10729_o;
  wire [31:0] n10730_o;
  wire [35:0] n10732_o;
  wire [35:0] n10733_o;
  wire [35:0] n10734_o;
  wire n10735_o;
  wire [37:0] n10737_o;
  wire [1:0] n10738_o;
  wire [1:0] n10739_o;
  wire [1:0] n10740_o;
  wire [35:0] n10741_o;
  wire [37:0] n10743_o;
  wire [37:0] n10744_o;
  wire [37:0] n10745_o;
  wire n10746_o;
  wire [38:0] n10748_o;
  wire [39:0] n10750_o;
  wire n10751_o;
  wire n10752_o;
  wire n10753_o;
  wire [38:0] n10754_o;
  wire [39:0] n10756_o;
  wire [39:0] n10757_o;
  wire [39:0] n10758_o;
  wire [39:0] n10759_o;
  wire [7:0] n10760_o;
  wire [7:0] n10761_o;
  wire [7:0] n10762_o;
  wire [31:0] n10763_o;
  wire n10764_o;
  wire n10765_o;
  wire [38:0] n10766_o;
  wire [39:0] n10767_o;
  wire [39:0] n10768_o;
  wire n10769_o;
  wire [1:0] n10770_o;
  wire [37:0] n10771_o;
  wire [39:0] n10772_o;
  wire [39:0] n10773_o;
  wire n10774_o;
  wire [3:0] n10775_o;
  wire [35:0] n10776_o;
  wire [39:0] n10777_o;
  wire [39:0] n10778_o;
  wire n10779_o;
  wire [7:0] n10780_o;
  wire [23:0] n10781_o;
  wire [31:0] n10782_o;
  wire [31:0] n10783_o;
  wire [31:0] n10784_o;
  wire n10785_o;
  wire [15:0] n10786_o;
  wire [15:0] n10787_o;
  wire [31:0] n10788_o;
  wire [31:0] n10789_o;
  wire [7:0] n10790_o;
  wire [31:0] n10791_o;
  wire [7:0] n10792_o;
  wire [39:0] n10793_o;
  localparam [39:0] n10794_o = 40'b0000000000000000000000000000000000000000;
  wire [39:0] n10796_o;
  localparam [39:0] n10798_o = 40'b1111111111111111111111111111111111111111;
  wire [39:0] n10800_o;
  wire [39:0] n10801_o;
  wire [39:0] n10802_o;
  wire n10803_o;
  wire n10804_o;
  wire n10805_o;
  wire n10806_o;
  wire n10807_o;
  wire n10808_o;
  wire n10809_o;
  wire n10810_o;
  wire n10811_o;
  wire n10812_o;
  wire n10820_o;
  wire n10821_o;
  wire n10822_o;
  wire n10823_o;
  wire n10824_o;
  wire n10825_o;
  wire n10826_o;
  wire n10827_o;
  wire n10828_o;
  wire n10829_o;
  wire n10837_o;
  wire n10838_o;
  wire n10839_o;
  wire n10840_o;
  wire n10841_o;
  wire n10842_o;
  wire n10843_o;
  wire n10844_o;
  wire n10845_o;
  wire n10846_o;
  wire n10854_o;
  wire n10855_o;
  wire n10856_o;
  wire n10857_o;
  wire n10858_o;
  wire n10859_o;
  wire n10860_o;
  wire n10861_o;
  wire n10862_o;
  wire n10863_o;
  wire n10871_o;
  wire n10872_o;
  wire n10873_o;
  wire n10874_o;
  wire n10875_o;
  wire n10876_o;
  wire n10877_o;
  wire n10878_o;
  wire n10879_o;
  wire n10880_o;
  wire n10888_o;
  wire n10889_o;
  wire n10890_o;
  wire n10891_o;
  wire n10892_o;
  wire n10893_o;
  wire n10894_o;
  wire n10895_o;
  wire n10896_o;
  wire n10897_o;
  wire n10905_o;
  wire n10906_o;
  wire n10907_o;
  wire n10908_o;
  wire n10909_o;
  wire n10910_o;
  wire n10911_o;
  wire n10912_o;
  wire n10913_o;
  wire n10914_o;
  wire n10922_o;
  wire n10923_o;
  wire n10924_o;
  wire n10925_o;
  wire n10926_o;
  wire n10927_o;
  wire n10928_o;
  wire n10929_o;
  wire n10930_o;
  wire n10931_o;
  wire n10939_o;
  wire n10940_o;
  wire n10941_o;
  wire n10942_o;
  wire n10943_o;
  wire n10944_o;
  wire n10945_o;
  wire n10946_o;
  wire n10947_o;
  wire n10948_o;
  wire n10956_o;
  wire n10957_o;
  wire n10958_o;
  wire n10959_o;
  wire n10960_o;
  wire n10961_o;
  wire n10962_o;
  wire n10963_o;
  wire n10964_o;
  wire n10965_o;
  wire n10973_o;
  wire n10974_o;
  wire n10975_o;
  wire n10976_o;
  wire n10977_o;
  wire n10978_o;
  wire n10979_o;
  wire n10980_o;
  wire n10981_o;
  wire n10982_o;
  wire n10990_o;
  wire n10991_o;
  wire n10992_o;
  wire n10993_o;
  wire n10994_o;
  wire n10995_o;
  wire n10996_o;
  wire n10997_o;
  wire n10998_o;
  wire n10999_o;
  wire n11007_o;
  wire n11008_o;
  wire n11009_o;
  wire n11010_o;
  wire n11011_o;
  wire n11012_o;
  wire n11013_o;
  wire n11014_o;
  wire n11015_o;
  wire n11016_o;
  wire n11024_o;
  wire n11025_o;
  wire n11026_o;
  wire n11027_o;
  wire n11028_o;
  wire n11029_o;
  wire n11030_o;
  wire n11031_o;
  wire n11032_o;
  wire n11033_o;
  wire n11041_o;
  wire n11042_o;
  wire n11043_o;
  wire n11044_o;
  wire n11045_o;
  wire n11046_o;
  wire n11047_o;
  wire n11048_o;
  wire n11049_o;
  wire n11050_o;
  wire n11058_o;
  wire n11059_o;
  wire n11060_o;
  wire n11061_o;
  wire n11062_o;
  wire n11063_o;
  wire n11064_o;
  wire n11065_o;
  wire n11066_o;
  wire n11067_o;
  wire n11075_o;
  wire n11076_o;
  wire n11077_o;
  wire n11078_o;
  wire n11079_o;
  wire n11080_o;
  wire n11081_o;
  wire n11082_o;
  wire n11083_o;
  wire n11084_o;
  wire n11092_o;
  wire n11093_o;
  wire n11094_o;
  wire n11095_o;
  wire n11096_o;
  wire n11097_o;
  wire n11098_o;
  wire n11099_o;
  wire n11100_o;
  wire n11101_o;
  wire n11109_o;
  wire n11110_o;
  wire n11111_o;
  wire n11112_o;
  wire n11113_o;
  wire n11114_o;
  wire n11115_o;
  wire n11116_o;
  wire n11117_o;
  wire n11118_o;
  wire n11126_o;
  wire n11127_o;
  wire n11128_o;
  wire n11129_o;
  wire n11130_o;
  wire n11131_o;
  wire n11132_o;
  wire n11133_o;
  wire n11134_o;
  wire n11135_o;
  wire n11143_o;
  wire n11144_o;
  wire n11145_o;
  wire n11146_o;
  wire n11147_o;
  wire n11148_o;
  wire n11149_o;
  wire n11150_o;
  wire n11151_o;
  wire n11152_o;
  wire n11160_o;
  wire n11161_o;
  wire n11162_o;
  wire n11163_o;
  wire n11164_o;
  wire n11165_o;
  wire n11166_o;
  wire n11167_o;
  wire n11168_o;
  wire n11169_o;
  wire n11177_o;
  wire n11178_o;
  wire n11179_o;
  wire n11180_o;
  wire n11181_o;
  wire n11182_o;
  wire n11183_o;
  wire n11184_o;
  wire n11185_o;
  wire n11186_o;
  wire n11194_o;
  wire n11195_o;
  wire n11196_o;
  wire n11197_o;
  wire n11198_o;
  wire n11199_o;
  wire n11200_o;
  wire n11201_o;
  wire n11202_o;
  wire n11203_o;
  wire n11211_o;
  wire n11212_o;
  wire n11213_o;
  wire n11214_o;
  wire n11215_o;
  wire n11216_o;
  wire n11217_o;
  wire n11218_o;
  wire n11219_o;
  wire n11220_o;
  wire n11228_o;
  wire n11229_o;
  wire n11230_o;
  wire n11231_o;
  wire n11232_o;
  wire n11233_o;
  wire n11234_o;
  wire n11235_o;
  wire n11236_o;
  wire n11237_o;
  wire n11245_o;
  wire n11246_o;
  wire n11247_o;
  wire n11248_o;
  wire n11249_o;
  wire n11250_o;
  wire n11251_o;
  wire n11252_o;
  wire n11253_o;
  wire n11254_o;
  wire n11262_o;
  wire n11263_o;
  wire n11264_o;
  wire n11265_o;
  wire n11266_o;
  wire n11267_o;
  wire n11268_o;
  wire n11269_o;
  wire n11270_o;
  wire n11271_o;
  wire n11279_o;
  wire n11280_o;
  wire n11281_o;
  wire n11282_o;
  wire n11283_o;
  wire n11284_o;
  wire n11285_o;
  wire n11286_o;
  wire n11287_o;
  wire n11288_o;
  wire n11296_o;
  wire n11297_o;
  wire n11298_o;
  wire n11299_o;
  wire n11300_o;
  wire n11301_o;
  wire n11302_o;
  wire n11303_o;
  wire n11304_o;
  wire n11305_o;
  wire n11313_o;
  wire n11314_o;
  wire n11315_o;
  wire n11316_o;
  wire n11317_o;
  wire n11318_o;
  wire n11319_o;
  wire n11320_o;
  wire n11321_o;
  wire n11322_o;
  wire n11330_o;
  wire n11331_o;
  wire n11332_o;
  wire n11333_o;
  wire n11334_o;
  wire n11335_o;
  wire n11336_o;
  wire n11337_o;
  wire n11338_o;
  wire n11339_o;
  wire n11347_o;
  wire n11348_o;
  wire n11349_o;
  wire n11350_o;
  wire n11351_o;
  wire n11352_o;
  wire n11353_o;
  wire n11354_o;
  wire n11355_o;
  wire n11356_o;
  wire n11364_o;
  wire n11365_o;
  wire n11366_o;
  wire n11367_o;
  wire n11368_o;
  wire n11369_o;
  wire n11370_o;
  wire n11371_o;
  wire n11372_o;
  wire n11373_o;
  wire n11381_o;
  wire n11382_o;
  wire n11383_o;
  wire n11384_o;
  wire n11385_o;
  wire n11386_o;
  wire n11387_o;
  wire n11388_o;
  wire n11389_o;
  wire n11390_o;
  wire n11398_o;
  wire n11399_o;
  wire n11400_o;
  wire n11401_o;
  wire n11402_o;
  wire n11403_o;
  wire n11404_o;
  wire n11405_o;
  wire n11406_o;
  wire n11407_o;
  wire n11415_o;
  wire n11416_o;
  wire n11417_o;
  wire n11418_o;
  wire n11419_o;
  wire n11420_o;
  wire n11421_o;
  wire n11422_o;
  wire n11423_o;
  wire n11424_o;
  wire n11432_o;
  wire n11433_o;
  wire n11434_o;
  wire n11435_o;
  wire n11436_o;
  wire n11437_o;
  wire n11438_o;
  wire n11439_o;
  wire n11440_o;
  wire n11441_o;
  wire n11449_o;
  wire n11450_o;
  wire n11451_o;
  wire n11452_o;
  wire n11453_o;
  wire n11454_o;
  wire n11455_o;
  wire n11456_o;
  wire n11457_o;
  wire n11458_o;
  wire n11459_o;
  wire n11460_o;
  wire n11461_o;
  wire n11462_o;
  wire n11463_o;
  wire n11464_o;
  wire n11465_o;
  wire n11466_o;
  wire n11467_o;
  wire n11468_o;
  wire [5:0] n11470_o;
  wire [5:0] n11471_o;
  wire [5:0] n11472_o;
  wire [3:0] n11473_o;
  wire n11475_o;
  wire [3:0] n11476_o;
  wire n11478_o;
  wire [3:0] n11479_o;
  wire n11481_o;
  wire [3:0] n11482_o;
  wire n11484_o;
  wire [3:0] n11486_o;
  wire n11488_o;
  wire [3:0] n11489_o;
  wire n11491_o;
  wire [3:0] n11493_o;
  wire n11495_o;
  wire [3:0] n11497_o;
  wire [3:0] n11498_o;
  wire [3:0] n11499_o;
  wire n11501_o;
  wire [3:0] n11502_o;
  wire [3:0] n11504_o;
  wire [1:0] n11505_o;
  wire n11506_o;
  wire n11507_o;
  wire n11508_o;
  wire n11510_o;
  wire [3:0] n11511_o;
  wire [3:0] n11512_o;
  wire [1:0] n11513_o;
  wire [1:0] n11515_o;
  wire [3:0] n11516_o;
  wire [3:0] n11519_o;
  wire [1:0] n11520_o;
  wire [2:0] n11521_o;
  wire [1:0] n11522_o;
  wire [1:0] n11523_o;
  wire n11524_o;
  wire n11526_o;
  wire [3:0] n11527_o;
  wire [3:0] n11529_o;
  wire [2:0] n11530_o;
  wire n11531_o;
  wire n11533_o;
  wire n11534_o;
  wire n11535_o;
  wire n11536_o;
  wire n11538_o;
  wire [3:0] n11539_o;
  wire [3:0] n11541_o;
  wire [2:0] n11542_o;
  wire n11543_o;
  wire n11544_o;
  wire [1:0] n11545_o;
  wire [1:0] n11547_o;
  wire [3:0] n11548_o;
  wire [3:0] n11549_o;
  wire [2:0] n11550_o;
  wire [2:0] n11552_o;
  localparam [4:0] n11553_o = 5'b11111;
  wire [1:0] n11555_o;
  wire n11557_o;
  wire n11559_o;
  wire n11560_o;
  wire n11562_o;
  wire n11563_o;
  wire n11566_o;
  wire n11567_o;
  wire n11568_o;
  wire n11570_o;
  wire n11571_o;
  wire n11572_o;
  wire n11574_o;
  wire n11575_o;
  wire [1:0] n11576_o;
  wire n11577_o;
  wire n11578_o;
  wire n11579_o;
  wire n11580_o;
  wire n11581_o;
  wire n11584_o;
  wire [1:0] n11589_o;
  wire n11590_o;
  wire n11592_o;
  wire n11593_o;
  wire n11595_o;
  wire n11597_o;
  wire n11598_o;
  wire n11599_o;
  wire n11601_o;
  wire [2:0] n11602_o;
  reg n11603_o;
  wire n11605_o;
  wire n11607_o;
  wire n11608_o;
  wire n11609_o;
  wire n11611_o;
  wire n11612_o;
  wire n11614_o;
  wire [3:0] n11615_o;
  reg n11618_o;
  reg n11620_o;
  wire n11621_o;
  wire n11622_o;
  wire n11624_o;
  wire n11625_o;
  wire n11627_o;
  wire n11628_o;
  wire [30:0] n11629_o;
  wire [31:0] n11630_o;
  wire n11631_o;
  wire n11632_o;
  wire [30:0] n11633_o;
  wire [31:0] n11634_o;
  wire [1:0] n11635_o;
  wire n11637_o;
  wire n11639_o;
  wire n11641_o;
  wire n11642_o;
  wire [1:0] n11643_o;
  wire n11644_o;
  reg n11645_o;
  wire n11646_o;
  reg n11647_o;
  wire [6:0] n11649_o;
  wire [15:0] n11650_o;
  wire [6:0] n11651_o;
  wire n11652_o;
  wire n11653_o;
  wire [31:0] n11654_o;
  wire [31:0] n11655_o;
  wire n11656_o;
  wire n11657_o;
  wire [31:0] n11658_o;
  wire n11663_o;
  wire [1:0] n11664_o;
  wire n11666_o;
  wire n11668_o;
  wire n11670_o;
  wire n11671_o;
  wire n11673_o;
  wire [2:0] n11674_o;
  reg [5:0] n11679_o;
  wire [1:0] n11680_o;
  wire n11682_o;
  wire n11684_o;
  wire n11686_o;
  wire n11687_o;
  wire n11689_o;
  wire [2:0] n11690_o;
  reg [5:0] n11695_o;
  wire [5:0] n11696_o;
  wire [1:0] n11698_o;
  wire n11700_o;
  wire n11701_o;
  wire n11702_o;
  wire n11703_o;
  wire n11704_o;
  wire [5:0] n11705_o;
  wire [2:0] n11706_o;
  wire [2:0] n11707_o;
  wire n11709_o;
  wire [2:0] n11712_o;
  wire [5:0] n11713_o;
  wire [5:0] n11714_o;
  wire [5:0] n11716_o;
  localparam [33:0] n11719_o = 34'b0000000000000000000000000000000000;
  wire n11723_o;
  wire [5:0] n11724_o;
  wire [5:0] n11726_o;
  wire [30:0] n11728_o;
  wire [31:0] n11730_o;
  wire [30:0] n11731_o;
  wire [31:0] n11733_o;
  wire [31:0] n11734_o;
  wire [32:0] n11735_o;
  wire [1:0] n11736_o;
  wire n11739_o;
  wire n11742_o;
  wire n11744_o;
  wire n11745_o;
  wire [1:0] n11746_o;
  wire n11747_o;
  reg n11748_o;
  wire n11749_o;
  reg n11750_o;
  wire [7:0] n11752_o;
  wire [15:0] n11753_o;
  wire [6:0] n11754_o;
  wire [31:0] n11755_o;
  wire [32:0] n11757_o;
  wire [32:0] n11758_o;
  wire n11760_o;
  wire n11761_o;
  wire n11762_o;
  wire n11763_o;
  wire n11764_o;
  wire n11766_o;
  wire n11768_o;
  wire n11769_o;
  wire n11770_o;
  wire [1:0] n11771_o;
  wire n11772_o;
  wire n11774_o;
  wire n11775_o;
  wire n11777_o;
  wire n11779_o;
  wire n11780_o;
  wire n11781_o;
  wire n11783_o;
  wire [2:0] n11784_o;
  reg n11785_o;
  wire n11786_o;
  wire n11788_o;
  wire n11789_o;
  wire [1:0] n11790_o;
  wire [7:0] n11791_o;
  wire [7:0] n11792_o;
  wire [7:0] n11793_o;
  wire n11794_o;
  wire n11796_o;
  wire [15:0] n11797_o;
  wire [15:0] n11798_o;
  wire [15:0] n11799_o;
  wire n11800_o;
  wire n11802_o;
  wire n11804_o;
  wire n11805_o;
  wire [31:0] n11806_o;
  wire [31:0] n11807_o;
  wire [31:0] n11808_o;
  wire n11809_o;
  wire n11811_o;
  wire [2:0] n11812_o;
  wire [7:0] n11813_o;
  wire [7:0] n11814_o;
  reg [7:0] n11816_o;
  wire [7:0] n11817_o;
  wire [7:0] n11818_o;
  reg [7:0] n11820_o;
  wire [15:0] n11821_o;
  reg [15:0] n11823_o;
  reg n11824_o;
  wire n11825_o;
  wire n11826_o;
  wire n11827_o;
  wire n11829_o;
  wire [1:0] n11830_o;
  wire [7:0] n11831_o;
  wire [7:0] n11832_o;
  wire [7:0] n11833_o;
  wire n11834_o;
  wire n11835_o;
  wire n11836_o;
  wire n11838_o;
  wire [15:0] n11839_o;
  wire [15:0] n11840_o;
  wire [15:0] n11841_o;
  wire n11842_o;
  wire n11843_o;
  wire n11844_o;
  wire n11846_o;
  wire n11848_o;
  wire n11849_o;
  wire [31:0] n11850_o;
  wire [31:0] n11851_o;
  wire [31:0] n11852_o;
  wire n11853_o;
  wire n11854_o;
  wire n11855_o;
  wire n11857_o;
  wire [2:0] n11858_o;
  wire [7:0] n11859_o;
  wire [7:0] n11860_o;
  reg [7:0] n11862_o;
  wire [7:0] n11863_o;
  wire [7:0] n11864_o;
  reg [7:0] n11866_o;
  wire [15:0] n11867_o;
  reg [15:0] n11869_o;
  reg n11870_o;
  wire n11871_o;
  wire n11872_o;
  wire [31:0] n11873_o;
  wire [31:0] n11874_o;
  wire [31:0] n11875_o;
  wire [31:0] n11876_o;
  wire [31:0] n11877_o;
  wire n11878_o;
  wire [31:0] n11879_o;
  wire [31:0] n11880_o;
  wire n11882_o;
  wire n11883_o;
  wire n11885_o;
  wire n11887_o;
  wire n11888_o;
  wire n11890_o;
  wire n11891_o;
  wire n11893_o;
  wire n11894_o;
  wire n11895_o;
  wire n11897_o;
  wire n11899_o;
  wire [5:0] n11901_o;
  wire n11903_o;
  wire [5:0] n11905_o;
  wire n11907_o;
  wire [5:0] n11909_o;
  wire n11911_o;
  wire [5:0] n11913_o;
  wire n11915_o;
  wire [5:0] n11917_o;
  wire n11919_o;
  wire [5:0] n11921_o;
  wire [5:0] n11922_o;
  wire [5:0] n11923_o;
  wire [5:0] n11924_o;
  wire [5:0] n11925_o;
  wire [5:0] n11926_o;
  wire [5:0] n11927_o;
  wire [5:0] n11929_o;
  wire n11931_o;
  wire n11933_o;
  wire [5:0] n11935_o;
  wire n11937_o;
  wire [5:0] n11939_o;
  wire n11941_o;
  wire [5:0] n11943_o;
  wire [5:0] n11944_o;
  wire [5:0] n11945_o;
  wire [5:0] n11946_o;
  wire n11948_o;
  wire n11950_o;
  wire [5:0] n11952_o;
  wire [5:0] n11953_o;
  wire n11955_o;
  wire [2:0] n11956_o;
  wire [5:0] n11958_o;
  wire n11960_o;
  wire [3:0] n11961_o;
  wire [5:0] n11963_o;
  wire n11965_o;
  wire [4:0] n11966_o;
  wire [5:0] n11968_o;
  wire n11970_o;
  wire [5:0] n11971_o;
  reg [5:0] n11973_o;
  wire n11974_o;
  wire n11975_o;
  wire [5:0] n11976_o;
  wire [5:0] n11977_o;
  wire n11978_o;
  wire n11979_o;
  wire n11980_o;
  wire n11981_o;
  wire [5:0] n11983_o;
  wire [5:0] n11984_o;
  wire n11985_o;
  wire n11986_o;
  wire n11987_o;
  wire [5:0] n11989_o;
  wire [5:0] n11990_o;
  wire [5:0] n11991_o;
  wire n11992_o;
  wire n11993_o;
  wire n11994_o;
  wire [5:0] n11996_o;
  wire [5:0] n11998_o;
  wire n12000_o;
  wire [5:0] n12001_o;
  wire n12002_o;
  wire [5:0] n12003_o;
  wire n12004_o;
  wire [31:0] n12005_o;
  wire [31:0] n12006_o;
  wire [31:0] n12007_o;
  localparam [32:0] n12008_o = 33'b000000000000000000000000000000000;
  wire n12009_o;
  wire n12011_o;
  wire n12012_o;
  wire n12013_o;
  wire n12014_o;
  wire n12015_o;
  wire [31:0] n12016_o;
  wire [31:0] n12017_o;
  wire n12018_o;
  wire n12020_o;
  wire n12022_o;
  wire [32:0] n12024_o;
  wire [1:0] n12025_o;
  wire n12026_o;
  localparam [23:0] n12027_o = 24'b000000000000000000000000;
  localparam [23:0] n12028_o = 24'b000000000000000000000000;
  wire n12030_o;
  wire n12031_o;
  wire n12032_o;
  wire n12033_o;
  wire [22:0] n12034_o;
  wire n12036_o;
  wire n12037_o;
  localparam [15:0] n12038_o = 16'b0000000000000000;
  wire n12041_o;
  wire n12042_o;
  wire n12043_o;
  wire n12044_o;
  wire [14:0] n12045_o;
  wire n12047_o;
  wire n12049_o;
  wire n12050_o;
  wire n12051_o;
  wire n12053_o;
  wire n12054_o;
  wire n12055_o;
  wire n12056_o;
  wire n12058_o;
  wire [2:0] n12059_o;
  wire n12060_o;
  reg n12061_o;
  wire [6:0] n12062_o;
  wire [6:0] n12063_o;
  reg [6:0] n12064_o;
  wire n12065_o;
  wire n12066_o;
  reg n12067_o;
  wire [14:0] n12068_o;
  wire [14:0] n12069_o;
  reg [14:0] n12070_o;
  wire n12071_o;
  reg n12072_o;
  wire [7:0] n12074_o;
  reg n12078_o;
  wire [7:0] n12079_o;
  wire [7:0] n12080_o;
  wire [7:0] n12081_o;
  wire [7:0] n12082_o;
  reg [7:0] n12083_o;
  wire [15:0] n12084_o;
  wire [15:0] n12085_o;
  wire [15:0] n12086_o;
  wire [15:0] n12087_o;
  reg [15:0] n12088_o;
  wire [7:0] n12092_o;
  wire [7:0] n12093_o;
  wire [7:0] n12094_o;
  wire [65:0] n12096_o;
  wire [30:0] n12097_o;
  wire [31:0] n12098_o;
  wire [65:0] n12099_o;
  wire n12103_o;
  wire [7:0] n12104_o;
  wire [7:0] n12105_o;
  wire n12106_o;
  wire [7:0] n12107_o;
  wire [7:0] n12108_o;
  wire n12109_o;
  wire [7:0] n12110_o;
  wire [7:0] n12111_o;
  wire [7:0] n12112_o;
  wire [7:0] n12113_o;
  wire [7:0] n12114_o;
  wire [7:0] n12115_o;
  wire n12116_o;
  wire n12117_o;
  wire n12118_o;
  wire n12119_o;
  wire [7:0] n12120_o;
  wire n12122_o;
  wire [7:0] n12124_o;
  wire n12126_o;
  wire [15:0] n12128_o;
  wire n12130_o;
  wire n12133_o;
  wire [1:0] n12134_o;
  wire [1:0] n12136_o;
  wire [2:0] n12137_o;
  wire [2:0] n12139_o;
  wire [2:0] n12141_o;
  wire n12144_o;
  wire n12145_o;
  wire n12146_o;
  wire [1:0] n12147_o;
  wire n12148_o;
  wire [2:0] n12149_o;
  wire n12150_o;
  wire [3:0] n12151_o;
  wire n12152_o;
  wire n12153_o;
  wire n12154_o;
  wire [1:0] n12155_o;
  wire [1:0] n12156_o;
  wire [1:0] n12157_o;
  wire [1:0] n12158_o;
  wire n12160_o;
  wire n12161_o;
  wire n12162_o;
  wire n12163_o;
  wire n12164_o;
  wire [1:0] n12165_o;
  wire n12166_o;
  wire [2:0] n12167_o;
  wire n12168_o;
  wire [3:0] n12169_o;
  wire n12170_o;
  wire n12171_o;
  wire [1:0] n12172_o;
  wire n12173_o;
  wire [2:0] n12174_o;
  wire n12175_o;
  wire [3:0] n12176_o;
  wire [3:0] n12177_o;
  wire [3:0] n12178_o;
  wire [3:0] n12179_o;
  wire n12181_o;
  wire n12182_o;
  wire n12185_o;
  wire n12188_o;
  wire n12189_o;
  wire n12190_o;
  wire n12191_o;
  wire n12192_o;
  wire n12193_o;
  wire n12195_o;
  wire n12196_o;
  wire n12198_o;
  wire n12199_o;
  wire n12200_o;
  wire n12201_o;
  wire n12202_o;
  wire [1:0] n12204_o;
  wire [3:0] n12206_o;
  wire [3:0] n12208_o;
  wire [3:0] n12209_o;
  wire [3:0] n12210_o;
  wire [3:0] n12211_o;
  wire [3:0] n12212_o;
  wire [3:0] n12213_o;
  wire [3:0] n12214_o;
  wire n12215_o;
  wire n12216_o;
  wire [3:0] n12217_o;
  wire n12218_o;
  wire n12219_o;
  wire n12220_o;
  wire n12222_o;
  wire n12223_o;
  wire n12224_o;
  wire n12225_o;
  wire n12226_o;
  wire n12227_o;
  wire n12228_o;
  wire n12229_o;
  wire n12230_o;
  wire n12231_o;
  wire n12232_o;
  wire n12233_o;
  wire n12234_o;
  wire n12235_o;
  wire n12236_o;
  wire n12237_o;
  wire n12238_o;
  wire n12239_o;
  wire n12241_o;
  wire n12243_o;
  wire n12245_o;
  wire n12246_o;
  wire n12247_o;
  wire [1:0] n12248_o;
  wire [3:0] n12250_o;
  wire n12251_o;
  wire n12252_o;
  wire [1:0] n12253_o;
  wire [3:0] n12255_o;
  wire [3:0] n12256_o;
  wire [3:0] n12257_o;
  wire n12258_o;
  wire n12260_o;
  wire n12261_o;
  wire n12262_o;
  wire n12263_o;
  wire n12264_o;
  wire n12267_o;
  wire n12269_o;
  wire n12270_o;
  wire n12271_o;
  wire n12273_o;
  wire n12274_o;
  wire n12275_o;
  wire n12276_o;
  wire n12277_o;
  wire n12278_o;
  wire n12279_o;
  wire n12280_o;
  wire n12281_o;
  wire n12282_o;
  wire n12283_o;
  wire n12284_o;
  wire n12285_o;
  wire n12286_o;
  wire n12288_o;
  wire n12289_o;
  wire n12292_o;
  wire n12293_o;
  wire n12294_o;
  wire n12295_o;
  wire n12296_o;
  wire [1:0] n12297_o;
  wire n12299_o;
  wire n12300_o;
  wire n12301_o;
  wire n12302_o;
  wire n12303_o;
  wire n12306_o;
  wire n12307_o;
  wire [1:0] n12308_o;
  wire n12309_o;
  wire n12310_o;
  wire n12311_o;
  wire n12312_o;
  wire n12313_o;
  wire n12314_o;
  wire n12315_o;
  wire n12316_o;
  wire n12317_o;
  wire n12318_o;
  wire n12319_o;
  wire n12320_o;
  wire n12321_o;
  wire n12322_o;
  wire n12323_o;
  wire n12324_o;
  wire n12325_o;
  wire n12326_o;
  wire n12327_o;
  wire n12328_o;
  wire n12329_o;
  wire n12330_o;
  wire n12332_o;
  wire n12333_o;
  wire n12334_o;
  wire n12335_o;
  wire n12336_o;
  wire n12337_o;
  wire n12339_o;
  wire n12340_o;
  wire n12341_o;
  wire n12342_o;
  wire [15:0] n12343_o;
  wire n12345_o;
  wire n12347_o;
  wire [15:0] n12348_o;
  wire n12350_o;
  wire n12351_o;
  wire n12352_o;
  wire n12355_o;
  wire [3:0] n12358_o;
  wire [3:0] n12359_o;
  wire [3:0] n12360_o;
  wire [3:0] n12361_o;
  wire [3:0] n12362_o;
  wire [3:0] n12363_o;
  wire [3:0] n12364_o;
  wire [3:0] n12365_o;
  wire [3:0] n12366_o;
  wire [1:0] n12367_o;
  wire [1:0] n12368_o;
  wire [1:0] n12369_o;
  wire [1:0] n12370_o;
  wire [1:0] n12371_o;
  wire [1:0] n12372_o;
  wire [1:0] n12373_o;
  wire n12374_o;
  wire n12375_o;
  wire n12376_o;
  wire n12377_o;
  wire n12378_o;
  wire n12379_o;
  wire n12380_o;
  wire n12381_o;
  wire n12382_o;
  wire [3:0] n12383_o;
  wire [3:0] n12384_o;
  wire [3:0] n12385_o;
  wire [3:0] n12386_o;
  wire [3:0] n12387_o;
  wire [3:0] n12388_o;
  wire [3:0] n12389_o;
  wire [3:0] n12390_o;
  wire [3:0] n12391_o;
  wire [3:0] n12392_o;
  wire [3:0] n12393_o;
  wire [3:0] n12394_o;
  wire [3:0] n12395_o;
  wire [4:0] n12396_o;
  wire [4:0] n12397_o;
  wire [4:0] n12398_o;
  wire [4:0] n12399_o;
  wire [4:0] n12400_o;
  wire [4:0] n12401_o;
  wire [4:0] n12402_o;
  wire [3:0] n12403_o;
  wire [3:0] n12404_o;
  wire [3:0] n12405_o;
  wire n12406_o;
  wire n12407_o;
  wire n12408_o;
  wire n12409_o;
  wire n12410_o;
  wire n12411_o;
  wire n12412_o;
  wire [3:0] n12413_o;
  wire [4:0] n12414_o;
  wire [4:0] n12415_o;
  wire [4:0] n12416_o;
  wire [2:0] n12417_o;
  wire [2:0] n12418_o;
  wire [2:0] n12419_o;
  wire [2:0] n12420_o;
  wire [2:0] n12421_o;
  wire [2:0] n12422_o;
  wire [2:0] n12423_o;
  wire [3:0] n12429_o;
  wire [7:0] n12430_o;
  wire [3:0] n12432_o;
  wire n12433_o;
  localparam [7:0] n12434_o = 8'b00000000;
  wire [3:0] n12436_o;
  wire n12437_o;
  wire [4:0] n12439_o;
  wire [4:0] n12440_o;
  wire [4:0] n12441_o;
  wire [4:0] n12442_o;
  wire [4:0] n12443_o;
  wire [7:0] n12444_o;
  wire n12451_o;
  wire n12452_o;
  wire n12453_o;
  wire n12454_o;
  wire n12456_o;
  wire n12457_o;
  wire n12458_o;
  wire n12461_o;
  wire [62:0] n12462_o;
  wire [63:0] n12463_o;
  wire n12464_o;
  wire [31:0] n12465_o;
  wire [32:0] n12466_o;
  wire [32:0] n12467_o;
  wire [32:0] n12468_o;
  wire [31:0] n12469_o;
  wire [32:0] n12470_o;
  wire [32:0] n12471_o;
  wire [32:0] n12472_o;
  wire [32:0] n12473_o;
  wire [32:0] n12474_o;
  wire [32:0] n12475_o;
  wire [30:0] n12476_o;
  wire n12477_o;
  wire n12479_o;
  wire [15:0] n12480_o;
  wire [31:0] n12482_o;
  wire [31:0] n12483_o;
  wire [31:0] n12484_o;
  wire n12486_o;
  wire n12487_o;
  wire n12488_o;
  wire n12489_o;
  wire n12490_o;
  wire n12491_o;
  wire [31:0] n12492_o;
  wire n12494_o;
  wire n12495_o;
  wire n12496_o;
  wire n12497_o;
  wire n12498_o;
  wire n12501_o;
  wire n12507_o;
  wire n12509_o;
  wire n12510_o;
  wire n12511_o;
  wire n12512_o;
  wire n12513_o;
  wire n12514_o;
  wire n12515_o;
  wire n12516_o;
  wire n12517_o;
  wire [31:0] n12519_o;
  wire [31:0] n12520_o;
  wire n12523_o;
  wire n12524_o;
  wire n12525_o;
  wire [63:0] n12526_o;
  wire [63:0] n12527_o;
  wire [63:0] n12528_o;
  wire [63:0] n12529_o;
  wire n12532_o;
  wire n12538_o;
  wire n12539_o;
  wire n12540_o;
  wire n12541_o;
  wire n12542_o;
  wire n12543_o;
  wire n12544_o;
  wire n12545_o;
  wire n12547_o;
  wire n12548_o;
  wire n12549_o;
  wire n12550_o;
  wire n12551_o;
  wire n12552_o;
  wire n12553_o;
  wire n12554_o;
  wire n12555_o;
  wire n12556_o;
  wire n12557_o;
  wire n12558_o;
  wire n12559_o;
  wire n12560_o;
  wire n12561_o;
  wire n12562_o;
  wire n12563_o;
  wire n12564_o;
  wire n12565_o;
  wire n12566_o;
  wire n12567_o;
  wire n12568_o;
  wire n12569_o;
  wire n12570_o;
  wire n12571_o;
  wire n12572_o;
  wire n12573_o;
  wire n12574_o;
  wire n12575_o;
  wire n12576_o;
  wire n12577_o;
  wire n12578_o;
  wire n12579_o;
  wire n12580_o;
  wire n12581_o;
  wire n12582_o;
  wire n12583_o;
  wire n12584_o;
  wire n12585_o;
  wire n12586_o;
  wire n12587_o;
  wire n12588_o;
  wire n12589_o;
  wire n12590_o;
  wire n12591_o;
  wire n12592_o;
  wire n12593_o;
  wire n12594_o;
  wire n12595_o;
  wire n12596_o;
  wire n12597_o;
  wire n12598_o;
  wire n12599_o;
  wire n12600_o;
  wire n12601_o;
  wire n12602_o;
  wire n12603_o;
  wire n12604_o;
  wire n12605_o;
  wire n12606_o;
  wire n12607_o;
  wire n12608_o;
  wire n12609_o;
  wire n12610_o;
  wire [3:0] n12611_o;
  wire [3:0] n12612_o;
  wire [3:0] n12613_o;
  wire [3:0] n12614_o;
  wire [3:0] n12615_o;
  wire [3:0] n12616_o;
  wire [3:0] n12617_o;
  wire [3:0] n12618_o;
  wire [15:0] n12619_o;
  wire [15:0] n12620_o;
  wire [31:0] n12621_o;
  wire n12622_o;
  wire n12624_o;
  wire n12625_o;
  wire n12626_o;
  wire n12627_o;
  wire n12628_o;
  wire [31:0] n12629_o;
  wire n12630_o;
  wire n12631_o;
  wire [63:0] n12632_o;
  wire [15:0] n12633_o;
  wire [15:0] n12634_o;
  wire [31:0] n12635_o;
  wire [31:0] n12636_o;
  wire [15:0] n12637_o;
  wire [15:0] n12638_o;
  wire [15:0] n12639_o;
  wire n12641_o;
  wire n12642_o;
  wire n12643_o;
  wire [15:0] n12644_o;
  wire [15:0] n12646_o;
  wire n12647_o;
  wire n12648_o;
  wire [32:0] n12649_o;
  wire [32:0] n12651_o;
  wire [32:0] n12652_o;
  wire [32:0] n12653_o;
  wire [16:0] n12655_o;
  wire [15:0] n12656_o;
  wire [32:0] n12657_o;
  wire [32:0] n12658_o;
  wire [32:0] n12659_o;
  wire n12660_o;
  wire [31:0] n12661_o;
  wire [31:0] n12662_o;
  wire [31:0] n12663_o;
  wire [30:0] n12664_o;
  wire n12665_o;
  wire [31:0] n12666_o;
  wire [31:0] n12667_o;
  wire [31:0] n12669_o;
  wire [31:0] n12670_o;
  wire [31:0] n12671_o;
  wire n12672_o;
  wire n12673_o;
  wire n12674_o;
  wire n12675_o;
  wire n12676_o;
  wire n12677_o;
  wire n12678_o;
  wire n12679_o;
  wire n12680_o;
  wire n12681_o;
  wire n12682_o;
  wire n12683_o;
  wire n12685_o;
  wire n12688_o;
  wire n12694_o;
  wire n12697_o;
  wire n12698_o;
  wire n12699_o;
  wire [63:0] n12701_o;
  wire [63:0] n12702_o;
  wire n12705_o;
  wire n12706_o;
  wire n12707_o;
  wire [63:0] n12708_o;
  wire n12710_o;
  wire n12713_o;
  wire n12714_o;
  wire n12715_o;
  wire n12716_o;
  wire [31:0] n12717_o;
  wire [32:0] n12719_o;
  wire [16:0] n12721_o;
  wire [15:0] n12722_o;
  wire [32:0] n12723_o;
  wire [32:0] n12724_o;
  wire n12727_o;
  wire n12728_o;
  wire [31:0] n12729_o;
  wire [31:0] n12731_o;
  wire [31:0] n12732_o;
  wire [31:0] n12733_o;
  wire [63:0] n12734_o;
  wire n12736_o;
  wire n12737_o;
  wire n12739_o;
  wire n12740_o;
  wire n12743_o;
  wire [31:0] n12753_o;
  wire [2:0] n12754_o;
  wire [3:0] n12755_o;
  reg [3:0] n12756_q;
  wire [8:0] n12757_o;
  wire [127:0] n12759_o;
  wire [63:0] n12760_o;
  reg [63:0] n12761_q;
  wire n12762_o;
  reg n12763_q;
  reg n12764_q;
  wire n12766_o;
  reg n12767_q;
  wire n12768_o;
  reg n12769_q;
  wire [63:0] n12771_o;
  reg [63:0] n12772_q;
  wire n12773_o;
  reg n12774_q;
  wire [63:0] n12776_o;
  reg [63:0] n12777_q;
  wire [63:0] n12778_o;
  wire n12780_o;
  reg n12781_q;
  wire [32:0] n12782_o;
  reg [32:0] n12783_q;
  wire n12784_o;
  reg n12785_q;
  wire [63:0] n12786_o;
  wire n12787_o;
  reg n12788_q;
  wire n12789_o;
  reg n12790_q;
  wire [31:0] n12793_o;
  wire [39:0] n12795_o;
  wire [31:0] n12796_o;
  wire [39:0] n12798_o;
  wire [4:0] n12799_o;
  wire n12800_o;
  reg n12801_q;
  wire n12802_o;
  reg n12803_q;
  wire n12804_o;
  reg n12805_q;
  wire n12806_o;
  reg n12807_q;
  wire n12808_o;
  reg n12809_q;
  wire n12810_o;
  reg n12811_q;
  wire n12812_o;
  reg n12813_q;
  wire [32:0] n12815_o;
  wire [32:0] n12816_o;
  wire [32:0] n12817_o;
  wire [31:0] n12818_o;
  wire [7:0] n12819_o;
  reg [7:0] n12820_q;
  reg [7:0] n12821_q;
  wire n12822_o;
  wire n12823_o;
  wire n12824_o;
  wire n12825_o;
  wire n12826_o;
  wire n12827_o;
  wire n12828_o;
  wire n12829_o;
  wire n12830_o;
  wire n12831_o;
  wire n12832_o;
  wire n12833_o;
  wire n12834_o;
  wire n12835_o;
  wire n12836_o;
  wire n12837_o;
  wire n12838_o;
  wire n12839_o;
  wire n12840_o;
  wire n12841_o;
  wire n12842_o;
  wire n12843_o;
  wire n12844_o;
  wire n12845_o;
  wire n12846_o;
  wire n12847_o;
  wire n12848_o;
  wire n12849_o;
  wire n12850_o;
  wire n12851_o;
  wire n12852_o;
  wire n12853_o;
  wire [1:0] n12854_o;
  reg n12855_o;
  wire [1:0] n12856_o;
  reg n12857_o;
  wire [1:0] n12858_o;
  reg n12859_o;
  wire [1:0] n12860_o;
  reg n12861_o;
  wire [1:0] n12862_o;
  reg n12863_o;
  wire [1:0] n12864_o;
  reg n12865_o;
  wire [1:0] n12866_o;
  reg n12867_o;
  wire [1:0] n12868_o;
  reg n12869_o;
  wire [1:0] n12870_o;
  reg n12871_o;
  wire [1:0] n12872_o;
  reg n12873_o;
  wire n12874_o;
  wire n12875_o;
  wire n12876_o;
  wire n12877_o;
  wire n12878_o;
  wire n12879_o;
  wire n12880_o;
  wire n12881_o;
  wire n12882_o;
  wire n12883_o;
  wire n12884_o;
  wire n12885_o;
  wire n12886_o;
  wire n12887_o;
  wire n12888_o;
  wire n12889_o;
  wire n12890_o;
  wire n12891_o;
  wire n12892_o;
  wire n12893_o;
  wire n12894_o;
  wire n12895_o;
  wire n12896_o;
  wire n12897_o;
  wire n12898_o;
  wire n12899_o;
  wire n12900_o;
  wire n12901_o;
  wire n12902_o;
  wire n12903_o;
  wire n12904_o;
  wire n12905_o;
  wire n12906_o;
  wire n12907_o;
  wire n12908_o;
  wire n12909_o;
  wire n12910_o;
  wire n12911_o;
  wire n12912_o;
  wire n12913_o;
  wire n12914_o;
  wire n12915_o;
  wire n12916_o;
  wire n12917_o;
  wire n12918_o;
  wire n12919_o;
  wire n12920_o;
  wire n12921_o;
  wire n12922_o;
  wire n12923_o;
  wire n12924_o;
  wire n12925_o;
  wire n12926_o;
  wire n12927_o;
  wire n12928_o;
  wire n12929_o;
  wire n12930_o;
  wire n12931_o;
  wire n12932_o;
  wire n12933_o;
  wire n12934_o;
  wire n12935_o;
  wire n12936_o;
  wire n12937_o;
  wire n12938_o;
  wire n12939_o;
  wire n12940_o;
  wire n12941_o;
  wire n12942_o;
  wire n12943_o;
  wire n12944_o;
  wire n12945_o;
  wire n12946_o;
  wire n12947_o;
  wire n12948_o;
  wire n12949_o;
  wire n12950_o;
  wire n12951_o;
  wire n12952_o;
  wire n12953_o;
  wire n12954_o;
  wire n12955_o;
  wire n12956_o;
  wire n12957_o;
  wire n12958_o;
  wire n12959_o;
  wire n12960_o;
  wire n12961_o;
  wire n12962_o;
  wire n12963_o;
  wire n12964_o;
  wire n12965_o;
  wire n12966_o;
  wire n12967_o;
  wire n12968_o;
  wire n12969_o;
  wire n12970_o;
  wire n12971_o;
  wire n12972_o;
  wire n12973_o;
  wire n12974_o;
  wire n12975_o;
  wire n12976_o;
  wire n12977_o;
  wire n12978_o;
  wire n12979_o;
  wire n12980_o;
  wire n12981_o;
  wire n12982_o;
  wire n12983_o;
  wire n12984_o;
  wire n12985_o;
  wire n12986_o;
  wire n12987_o;
  wire n12988_o;
  wire n12989_o;
  wire n12990_o;
  wire n12991_o;
  wire n12992_o;
  wire n12993_o;
  wire n12994_o;
  wire n12995_o;
  wire n12996_o;
  wire n12997_o;
  wire n12998_o;
  wire n12999_o;
  wire n13000_o;
  wire n13001_o;
  wire n13002_o;
  wire n13003_o;
  wire n13004_o;
  wire n13005_o;
  wire n13006_o;
  wire n13007_o;
  wire n13008_o;
  wire n13009_o;
  wire [31:0] n13010_o;
  wire n13011_o;
  wire n13012_o;
  wire n13013_o;
  wire n13014_o;
  wire n13015_o;
  wire n13016_o;
  wire n13017_o;
  wire n13018_o;
  wire n13019_o;
  wire n13020_o;
  wire n13021_o;
  wire n13022_o;
  wire n13023_o;
  wire n13024_o;
  wire n13025_o;
  wire n13026_o;
  wire n13027_o;
  wire n13028_o;
  wire n13029_o;
  wire n13030_o;
  wire n13031_o;
  wire n13032_o;
  wire n13033_o;
  wire n13034_o;
  wire n13035_o;
  wire n13036_o;
  wire n13037_o;
  wire n13038_o;
  wire n13039_o;
  wire n13040_o;
  wire n13041_o;
  wire n13042_o;
  wire [1:0] n13043_o;
  reg n13044_o;
  wire [1:0] n13045_o;
  reg n13046_o;
  wire [1:0] n13047_o;
  reg n13048_o;
  wire [1:0] n13049_o;
  reg n13050_o;
  wire [1:0] n13051_o;
  reg n13052_o;
  wire [1:0] n13053_o;
  reg n13054_o;
  wire [1:0] n13055_o;
  reg n13056_o;
  wire [1:0] n13057_o;
  reg n13058_o;
  wire [1:0] n13059_o;
  reg n13060_o;
  wire [1:0] n13061_o;
  reg n13062_o;
  wire n13063_o;
  wire n13064_o;
  wire n13065_o;
  wire n13066_o;
  wire n13067_o;
  wire n13068_o;
  wire n13069_o;
  wire n13070_o;
  wire n13071_o;
  wire n13072_o;
  wire n13073_o;
  wire n13074_o;
  wire n13075_o;
  wire n13076_o;
  wire n13077_o;
  wire n13078_o;
  wire n13079_o;
  wire n13080_o;
  wire n13081_o;
  wire n13082_o;
  wire n13083_o;
  wire n13084_o;
  wire n13085_o;
  wire n13086_o;
  wire n13087_o;
  wire n13088_o;
  wire n13089_o;
  wire n13090_o;
  wire n13091_o;
  wire n13092_o;
  wire n13093_o;
  wire n13094_o;
  wire n13095_o;
  wire n13096_o;
  wire n13097_o;
  wire n13098_o;
  wire n13099_o;
  wire n13100_o;
  wire n13101_o;
  wire n13102_o;
  wire n13103_o;
  wire n13104_o;
  wire n13105_o;
  wire n13106_o;
  wire n13107_o;
  wire n13108_o;
  wire n13109_o;
  wire n13110_o;
  wire n13111_o;
  wire n13112_o;
  wire n13113_o;
  wire n13114_o;
  wire n13115_o;
  wire n13116_o;
  wire n13117_o;
  wire n13118_o;
  wire n13119_o;
  wire n13120_o;
  wire n13121_o;
  wire n13122_o;
  wire n13123_o;
  wire n13124_o;
  wire n13125_o;
  wire n13126_o;
  wire n13127_o;
  wire n13128_o;
  wire n13129_o;
  wire n13130_o;
  wire n13131_o;
  wire n13132_o;
  wire n13133_o;
  wire n13134_o;
  wire n13135_o;
  wire n13136_o;
  wire n13137_o;
  wire n13138_o;
  wire n13139_o;
  wire n13140_o;
  wire n13141_o;
  wire n13142_o;
  wire n13143_o;
  wire n13144_o;
  wire n13145_o;
  wire n13146_o;
  wire n13147_o;
  wire n13148_o;
  wire n13149_o;
  wire n13150_o;
  wire n13151_o;
  wire n13152_o;
  wire n13153_o;
  wire n13154_o;
  wire n13155_o;
  wire n13156_o;
  wire n13157_o;
  wire n13158_o;
  wire n13159_o;
  wire n13160_o;
  wire n13161_o;
  wire n13162_o;
  wire n13163_o;
  wire n13164_o;
  wire n13165_o;
  wire n13166_o;
  wire n13167_o;
  wire n13168_o;
  wire n13169_o;
  wire n13170_o;
  wire n13171_o;
  wire n13172_o;
  wire n13173_o;
  wire n13174_o;
  wire n13175_o;
  wire n13176_o;
  wire n13177_o;
  wire n13178_o;
  wire n13179_o;
  wire n13180_o;
  wire n13181_o;
  wire n13182_o;
  wire n13183_o;
  wire n13184_o;
  wire n13185_o;
  wire n13186_o;
  wire n13187_o;
  wire n13188_o;
  wire n13189_o;
  wire n13190_o;
  wire n13191_o;
  wire n13192_o;
  wire n13193_o;
  wire n13194_o;
  wire n13195_o;
  wire n13196_o;
  wire n13197_o;
  wire n13198_o;
  wire n13199_o;
  wire n13200_o;
  wire n13201_o;
  wire n13202_o;
  wire n13203_o;
  wire n13204_o;
  wire n13205_o;
  wire n13206_o;
  wire n13207_o;
  wire n13208_o;
  wire n13209_o;
  wire n13210_o;
  wire n13211_o;
  wire n13212_o;
  wire [33:0] n13213_o;
  assign bf_ext_out = n12820_q;
  assign set_v_flag = n12688_o;
  assign flags = n12821_q;
  assign c_out = n10046_o;
  assign addsub_q = n10024_o;
  assign aluout = n9804_o;
  /* TG68K_ALU.vhd:86:16  */
  assign op1in = n12753_o; // (signal)
  /* TG68K_ALU.vhd:87:16  */
  assign addsub_a = n9912_o; // (signal)
  /* TG68K_ALU.vhd:88:16  */
  assign addsub_b = n9995_o; // (signal)
  /* TG68K_ALU.vhd:89:16  */
  assign notaddsub_b = n10007_o; // (signal)
  /* TG68K_ALU.vhd:90:16  */
  assign add_result = n10012_o; // (signal)
  /* TG68K_ALU.vhd:91:16  */
  assign addsub_ofl = n12754_o; // (signal)
  /* TG68K_ALU.vhd:92:16  */
  assign opaddsub = n9974_o; // (signal)
  /* TG68K_ALU.vhd:93:16  */
  assign c_in = n12755_o; // (signal)
  /* TG68K_ALU.vhd:94:16  */
  assign flag_z = n12141_o; // (signal)
  /* TG68K_ALU.vhd:95:16  */
  assign set_flags = n12179_o; // (signal)
  /* TG68K_ALU.vhd:96:16  */
  assign ccrin = n12115_o; // (signal)
  /* TG68K_ALU.vhd:97:16  */
  assign last_flags1 = n12756_q; // (signal)
  /* TG68K_ALU.vhd:100:16  */
  assign bcd_pur = n10052_o; // (signal)
  /* TG68K_ALU.vhd:101:16  */
  assign bcd_kor = n12757_o; // (signal)
  /* TG68K_ALU.vhd:102:16  */
  assign halve_carry = n10057_o; // (signal)
  /* TG68K_ALU.vhd:103:16  */
  assign vflag_a = n10110_o; // (signal)
  /* TG68K_ALU.vhd:104:16  */
  assign bcd_a_carry = n10113_o; // (signal)
  /* TG68K_ALU.vhd:105:16  */
  assign bcd_a = n10107_o; // (signal)
  /* TG68K_ALU.vhd:106:16  */
  assign result_mulu = n12759_o; // (signal)
  /* TG68K_ALU.vhd:107:16  */
  assign result_div = n12761_q; // (signal)
  /* TG68K_ALU.vhd:108:16  */
  assign result_div_pre = n12671_o; // (signal)
  /* TG68K_ALU.vhd:109:16  */
  assign set_mv_flag = n12501_o; // (signal)
  /* TG68K_ALU.vhd:110:16  */
  assign v_flag = n12763_q; // (signal)
  /* TG68K_ALU.vhd:112:16  */
  assign rot_rot = n11603_o; // (signal)
  /* TG68K_ALU.vhd:113:16  */
  assign rot_lsb = n11618_o; // (signal)
  /* TG68K_ALU.vhd:114:16  */
  assign rot_msb = n11620_o; // (signal)
  /* TG68K_ALU.vhd:115:16  */
  assign rot_x = n11656_o; // (signal)
  /* TG68K_ALU.vhd:116:16  */
  assign rot_c = n11657_o; // (signal)
  /* TG68K_ALU.vhd:117:16  */
  assign rot_out = n11658_o; // (signal)
  /* TG68K_ALU.vhd:118:16  */
  assign asl_vflag = n12764_q; // (signal)
  /* TG68K_ALU.vhd:120:16  */
  assign bit_number = n10154_o; // (signal)
  /* TG68K_ALU.vhd:121:16  */
  assign bits_out = n13010_o; // (signal)
  /* TG68K_ALU.vhd:122:16  */
  assign one_bit_in = n12875_o; // (signal)
  /* TG68K_ALU.vhd:123:16  */
  assign bchg = n12767_q; // (signal)
  /* TG68K_ALU.vhd:124:16  */
  assign bset = n12769_q; // (signal)
  /* TG68K_ALU.vhd:126:16  */
  assign mulu_sign = n12461_o; // (signal)
  /* TG68K_ALU.vhd:128:16  */
  assign muls_msb = n12456_o; // (signal)
  /* TG68K_ALU.vhd:129:16  */
  assign mulu_reg = n12772_q; // (signal)
  /* TG68K_ALU.vhd:130:16  */
  assign fasign = n12774_q; // (signal)
  /* TG68K_ALU.vhd:132:16  */
  assign faktorb = n12483_o; // (signal)
  /* TG68K_ALU.vhd:134:16  */
  assign div_reg = n12777_q; // (signal)
  /* TG68K_ALU.vhd:135:16  */
  assign div_quot = n12778_o; // (signal)
  /* TG68K_ALU.vhd:137:16  */
  assign div_neg = n12781_q; // (signal)
  /* TG68K_ALU.vhd:138:16  */
  assign div_bit = n12660_o; // (signal)
  /* TG68K_ALU.vhd:139:16  */
  assign div_sub = n12659_o; // (signal)
  /* TG68K_ALU.vhd:140:16  */
  assign div_over = n12783_q; // (signal)
  /* TG68K_ALU.vhd:141:16  */
  assign nozero = n12785_q; // (signal)
  /* TG68K_ALU.vhd:142:16  */
  assign div_qsign = n12631_o; // (signal)
  /* TG68K_ALU.vhd:143:16  */
  assign dividend = n12786_o; // (signal)
  /* TG68K_ALU.vhd:144:16  */
  assign divs = n12545_o; // (signal)
  /* TG68K_ALU.vhd:145:16  */
  assign signedop = n12788_q; // (signal)
  /* TG68K_ALU.vhd:146:16  */
  assign op1_sign = n12790_q; // (signal)
  /* TG68K_ALU.vhd:148:16  */
  assign op2outext = n12646_o; // (signal)
  /* TG68K_ALU.vhd:151:16  */
  assign datareg = n12793_o; // (signal)
  /* TG68K_ALU.vhd:153:16  */
  assign bf_datareg = n10713_o; // (signal)
  /* TG68K_ALU.vhd:154:16  */
  assign result = n12795_o; // (signal)
  /* TG68K_ALU.vhd:155:16  */
  assign result_tmp = n10802_o; // (signal)
  /* TG68K_ALU.vhd:156:16  */
  assign unshifted_bitmask = n12796_o; // (signal)
  /* TG68K_ALU.vhd:158:16  */
  assign inmux0 = n10768_o; // (signal)
  /* TG68K_ALU.vhd:159:16  */
  assign inmux1 = n10773_o; // (signal)
  /* TG68K_ALU.vhd:160:16  */
  assign inmux2 = n10778_o; // (signal)
  /* TG68K_ALU.vhd:161:16  */
  assign inmux3 = n10784_o; // (signal)
  /* TG68K_ALU.vhd:162:16  */
  assign shifted_bitmask = n10758_o; // (signal)
  /* TG68K_ALU.vhd:163:16  */
  assign bitmaskmux0 = n10745_o; // (signal)
  /* TG68K_ALU.vhd:164:16  */
  assign bitmaskmux1 = n10734_o; // (signal)
  /* TG68K_ALU.vhd:165:16  */
  assign bitmaskmux2 = n10723_o; // (signal)
  /* TG68K_ALU.vhd:166:16  */
  assign bitmaskmux3 = n10718_o; // (signal)
  /* TG68K_ALU.vhd:167:16  */
  assign bf_set2 = n10789_o; // (signal)
  /* TG68K_ALU.vhd:168:16  */
  assign shift = n12798_o; // (signal)
  /* TG68K_ALU.vhd:169:16  */
  assign bf_firstbit = n11472_o; // (signal)
  /* TG68K_ALU.vhd:170:16  */
  assign mux = n11549_o; // (signal)
  /* TG68K_ALU.vhd:171:16  */
  assign bitnr = n12799_o; // (signal)
  /* TG68K_ALU.vhd:172:16  */
  assign mask = datareg; // (signal)
  /* TG68K_ALU.vhd:173:16  */
  assign mask_not_zero = n11584_o; // (signal)
  /* TG68K_ALU.vhd:174:16  */
  assign bf_bset = n12801_q; // (signal)
  /* TG68K_ALU.vhd:175:16  */
  assign bf_nflag = n13064_o; // (signal)
  /* TG68K_ALU.vhd:176:16  */
  assign bf_bchg = n12803_q; // (signal)
  /* TG68K_ALU.vhd:177:16  */
  assign bf_ins = n12805_q; // (signal)
  /* TG68K_ALU.vhd:178:16  */
  assign bf_exts = n12807_q; // (signal)
  /* TG68K_ALU.vhd:179:16  */
  assign bf_fffo = n12809_q; // (signal)
  /* TG68K_ALU.vhd:180:16  */
  assign bf_d32 = n12811_q; // (signal)
  /* TG68K_ALU.vhd:181:16  */
  assign bf_s32 = n12813_q; // (signal)
  /* TG68K_ALU.vhd:187:16  */
  assign hot_msb = n13213_o; // (signal)
  /* TG68K_ALU.vhd:188:16  */
  assign vector = n12815_o; // (signal)
  /* TG68K_ALU.vhd:189:16  */
  assign result_bs = n12099_o; // (signal)
  /* TG68K_ALU.vhd:190:16  */
  assign bit_nr = n12003_o; // (signal)
  /* TG68K_ALU.vhd:191:16  */
  assign bit_msb = n11726_o; // (signal)
  /* TG68K_ALU.vhd:192:16  */
  assign bs_shift = n11716_o; // (signal)
  /* TG68K_ALU.vhd:193:16  */
  assign bs_shift_mod = n11973_o; // (signal)
  /* TG68K_ALU.vhd:194:16  */
  assign asl_over = n11758_o; // (signal)
  /* TG68K_ALU.vhd:195:16  */
  assign asl_over_xor = n12816_o; // (signal)
  /* TG68K_ALU.vhd:196:16  */
  assign asr_sign = n12817_o; // (signal)
  /* TG68K_ALU.vhd:197:16  */
  assign msb = n12078_o; // (signal)
  /* TG68K_ALU.vhd:198:16  */
  assign ring = n11696_o; // (signal)
  /* TG68K_ALU.vhd:199:16  */
  assign alu = n11880_o; // (signal)
  /* TG68K_ALU.vhd:200:16  */
  assign bsout = n12818_o; // (signal)
  /* TG68K_ALU.vhd:201:16  */
  assign bs_v = n11893_o; // (signal)
  /* TG68K_ALU.vhd:202:16  */
  assign bs_c = n12020_o; // (signal)
  /* TG68K_ALU.vhd:203:16  */
  assign bs_x = n11895_o; // (signal)
  /* TG68K_ALU.vhd:215:35  */
  assign n9794_o = op1in[7];
  /* TG68K_ALU.vhd:215:39  */
  assign n9795_o = n9794_o | exec_tas;
  assign n9796_o = op1in[31:8];
  assign n9797_o = op1in[6:0];
  /* TG68K_ALU.vhd:216:24  */
  assign n9798_o = exec[76];
  /* TG68K_ALU.vhd:217:41  */
  assign n9799_o = result[31:0];
  /* TG68K_ALU.vhd:219:57  */
  assign n9800_o = {26'b0, bf_firstbit};  //  uext
  /* TG68K_ALU.vhd:219:57  */
  assign n9801_o = bf_ffo_offset - n9800_o;
  /* TG68K_ALU.vhd:218:25  */
  assign n9802_o = bf_fffo ? n9801_o : n9799_o;
  assign n9803_o = {n9796_o, n9795_o, n9797_o};
  /* TG68K_ALU.vhd:216:17  */
  assign n9804_o = n9798_o ? n9802_o : n9803_o;
  /* TG68K_ALU.vhd:224:24  */
  assign n9805_o = exec[12];
  /* TG68K_ALU.vhd:224:45  */
  assign n9806_o = exec[13];
  /* TG68K_ALU.vhd:224:38  */
  assign n9807_o = n9805_o | n9806_o;
  /* TG68K_ALU.vhd:225:51  */
  assign n9808_o = bcd_a[7:0];
  /* TG68K_ALU.vhd:226:27  */
  assign n9809_o = exec[20];
  /* TG68K_ALU.vhd:226:41  */
  assign n9811_o = 1'b1 & n9809_o;
  /* TG68K_ALU.vhd:228:40  */
  assign n9812_o = exec[67];
  /* TG68K_ALU.vhd:228:60  */
  assign n9814_o = 1'b1 & n9812_o;
  /* TG68K_ALU.vhd:229:61  */
  assign n9815_o = result_mulu[31:0];
  /* TG68K_ALU.vhd:231:61  */
  assign n9816_o = result_mulu[63:32];
  /* TG68K_ALU.vhd:228:33  */
  assign n9817_o = n9814_o ? n9815_o : n9816_o;
  /* TG68K_ALU.vhd:241:27  */
  assign n9818_o = exec[21];
  /* TG68K_ALU.vhd:241:41  */
  assign n9820_o = 1'b1 & n9818_o;
  /* TG68K_ALU.vhd:242:38  */
  assign n9821_o = exe_opcode[15];
  /* TG68K_ALU.vhd:242:47  */
  assign n9823_o = n9821_o | 1'b0;
  /* TG68K_ALU.vhd:244:52  */
  assign n9824_o = result_div[47:32];
  /* TG68K_ALU.vhd:244:77  */
  assign n9825_o = result_div[15:0];
  /* TG68K_ALU.vhd:244:66  */
  assign n9826_o = {n9824_o, n9825_o};
  /* TG68K_ALU.vhd:246:40  */
  assign n9827_o = exec[68];
  /* TG68K_ALU.vhd:247:60  */
  assign n9828_o = result_div[63:32];
  /* TG68K_ALU.vhd:249:60  */
  assign n9829_o = result_div[31:0];
  /* TG68K_ALU.vhd:246:33  */
  assign n9830_o = n9827_o ? n9828_o : n9829_o;
  /* TG68K_ALU.vhd:242:25  */
  assign n9831_o = n9823_o ? n9826_o : n9830_o;
  /* TG68K_ALU.vhd:252:27  */
  assign n9832_o = exec[5];
  /* TG68K_ALU.vhd:253:41  */
  assign n9833_o = op2out | op1out;
  /* TG68K_ALU.vhd:254:27  */
  assign n9834_o = exec[6];
  /* TG68K_ALU.vhd:255:41  */
  assign n9835_o = op2out & op1out;
  /* TG68K_ALU.vhd:256:27  */
  assign n9836_o = exec[16];
  assign n9837_o = {exe_condition, exe_condition, exe_condition, exe_condition};
  assign n9838_o = {exe_condition, exe_condition, exe_condition, exe_condition};
  assign n9839_o = {n9837_o, n9838_o};
  /* TG68K_ALU.vhd:258:27  */
  assign n9840_o = exec[7];
  /* TG68K_ALU.vhd:259:41  */
  assign n9841_o = op2out ^ op1out;
  /* TG68K_ALU.vhd:261:27  */
  assign n9842_o = exec[85];
  /* TG68K_ALU.vhd:264:27  */
  assign n9843_o = exec[9];
  /* TG68K_ALU.vhd:266:27  */
  assign n9844_o = exec[81];
  /* TG68K_ALU.vhd:268:27  */
  assign n9845_o = exec[15];
  /* TG68K_ALU.vhd:269:40  */
  assign n9846_o = op1out[15:0];
  /* TG68K_ALU.vhd:269:61  */
  assign n9847_o = op1out[31:16];
  /* TG68K_ALU.vhd:269:53  */
  assign n9848_o = {n9846_o, n9847_o};
  /* TG68K_ALU.vhd:270:27  */
  assign n9849_o = exec[14];
  /* TG68K_ALU.vhd:272:27  */
  assign n9850_o = exec[75];
  /* TG68K_ALU.vhd:274:27  */
  assign n9851_o = exec[2];
  /* TG68K_ALU.vhd:276:38  */
  assign n9852_o = exe_opcode[9];
  /* TG68K_ALU.vhd:276:25  */
  assign n9854_o = n9852_o ? 8'b00000000 : flagssr;
  /* TG68K_ALU.vhd:281:27  */
  assign n9855_o = exec[77];
  /* TG68K_ALU.vhd:282:54  */
  assign n9856_o = n10024_o[11:8];
  /* TG68K_ALU.vhd:282:78  */
  assign n9857_o = n10024_o[3:0];
  /* TG68K_ALU.vhd:282:68  */
  assign n9858_o = {n9856_o, n9857_o};
  assign n9859_o = n10024_o[7:0];
  /* TG68K_ALU.vhd:281:17  */
  assign n9860_o = n9855_o ? n9858_o : n9859_o;
  assign n9861_o = {n9854_o, n12821_q};
  assign n9862_o = n9861_o[7:0];
  /* TG68K_ALU.vhd:274:17  */
  assign n9863_o = n9851_o ? n9862_o : n9860_o;
  assign n9864_o = n9861_o[15:8];
  assign n9865_o = n10024_o[15:8];
  /* TG68K_ALU.vhd:274:17  */
  assign n9866_o = n9851_o ? n9864_o : n9865_o;
  assign n9867_o = {n9866_o, n9863_o};
  /* TG68KdotC_Kernel.vhd:2260:130  */
  assign n9868_o = bf_datareg[15:0];
  /* TG68K_ALU.vhd:272:17  */
  assign n9869_o = n9850_o ? n9868_o : n9867_o;
  /* TG68KdotC_Kernel.vhd:2260:183  */
  assign n9870_o = bf_datareg[31:16];
  assign n9871_o = n10024_o[31:16];
  /* TG68K_ALU.vhd:272:17  */
  assign n9872_o = n9850_o ? n9870_o : n9871_o;
  /* TG68KdotC_Kernel.vhd:2260:153  */
  assign n9873_o = {n9872_o, n9869_o};
  /* TG68K_ALU.vhd:270:17  */
  assign n9874_o = n9849_o ? bits_out : n9873_o;
  /* TG68K_ALU.vhd:268:17  */
  assign n9875_o = n9845_o ? n9848_o : n9874_o;
  /* TG68K_ALU.vhd:266:17  */
  assign n9876_o = n9844_o ? bsout : n9875_o;
  /* TG68K_ALU.vhd:264:17  */
  assign n9877_o = n9843_o ? rot_out : n9876_o;
  /* TG68K_ALU.vhd:261:17  */
  assign n9878_o = n9842_o ? op2out : n9877_o;
  /* TG68K_ALU.vhd:258:17  */
  assign n9879_o = n9840_o ? n9841_o : n9878_o;
  /* TG68KdotC_Kernel.vhd:2260:94  */
  assign n9880_o = n9879_o[7:0];
  /* TG68K_ALU.vhd:256:17  */
  assign n9881_o = n9836_o ? n9839_o : n9880_o;
  /* TG68KdotC_Kernel.vhd:2260:82  */
  assign n9882_o = n9879_o[31:8];
  assign n9883_o = n10024_o[31:8];
  /* TG68K_ALU.vhd:256:17  */
  assign n9884_o = n9836_o ? n9883_o : n9882_o;
  assign n9885_o = {n9884_o, n9881_o};
  /* TG68K_ALU.vhd:254:17  */
  assign n9886_o = n9834_o ? n9835_o : n9885_o;
  /* TG68K_ALU.vhd:252:17  */
  assign n9887_o = n9832_o ? n9833_o : n9886_o;
  /* TG68K_ALU.vhd:241:17  */
  assign n9888_o = n9820_o ? n9831_o : n9887_o;
  /* TG68K_ALU.vhd:226:17  */
  assign n9889_o = n9811_o ? n9817_o : n9888_o;
  assign n9890_o = n9889_o[7:0];
  /* TG68K_ALU.vhd:224:17  */
  assign n9891_o = n9807_o ? n9808_o : n9890_o;
  assign n9892_o = n9889_o[31:8];
  assign n9893_o = n10024_o[31:8];
  /* TG68K_ALU.vhd:224:17  */
  assign n9894_o = n9807_o ? n9893_o : n9892_o;
  /* TG68K_ALU.vhd:293:24  */
  assign n9899_o = exec[29];
  /* TG68K_ALU.vhd:294:34  */
  assign n9900_o = sndopc[11];
  /* TG68K_ALU.vhd:295:51  */
  assign n9901_o = op1out[31];
  /* TG68K_ALU.vhd:295:62  */
  assign n9902_o = op1out[31];
  /* TG68K_ALU.vhd:295:55  */
  assign n9903_o = {n9901_o, n9902_o};
  /* TG68K_ALU.vhd:295:73  */
  assign n9904_o = op1out[31];
  /* TG68K_ALU.vhd:295:66  */
  assign n9905_o = {n9903_o, n9904_o};
  /* TG68K_ALU.vhd:295:84  */
  assign n9906_o = op1out[31:3];
  /* TG68K_ALU.vhd:295:77  */
  assign n9907_o = {n9905_o, n9906_o};
  /* TG68K_ALU.vhd:297:84  */
  assign n9908_o = sndopc[10:9];
  /* TG68K_ALU.vhd:297:77  */
  assign n9910_o = {30'b000000000000000000000000000000, n9908_o};
  /* TG68K_ALU.vhd:294:25  */
  assign n9911_o = n9900_o ? n9907_o : n9910_o;
  /* TG68K_ALU.vhd:293:17  */
  assign n9912_o = n9899_o ? n9911_o : op1out;
  /* TG68K_ALU.vhd:301:24  */
  assign n9913_o = exec[48];
  /* TG68K_ALU.vhd:301:17  */
  assign n9916_o = n9913_o ? 1'b1 : 1'b0;
  /* TG68K_ALU.vhd:309:24  */
  assign n9918_o = exec[78];
  /* TG68K_ALU.vhd:310:65  */
  assign n9919_o = op2out[7:4];
  /* TG68K_ALU.vhd:310:57  */
  assign n9921_o = {4'b0000, n9919_o};
  /* TG68K_ALU.vhd:310:78  */
  assign n9923_o = {n9921_o, 4'b0000};
  /* TG68K_ALU.vhd:310:95  */
  assign n9924_o = op2out[3:0];
  /* TG68K_ALU.vhd:310:87  */
  assign n9925_o = {n9923_o, n9924_o};
  /* TG68K_ALU.vhd:311:30  */
  assign n9926_o = ~execopc;
  /* TG68K_ALU.vhd:311:43  */
  assign n9927_o = exec[53];
  /* TG68K_ALU.vhd:311:55  */
  assign n9928_o = ~n9927_o;
  /* TG68K_ALU.vhd:311:35  */
  assign n9929_o = n9928_o & n9926_o;
  /* TG68K_ALU.vhd:311:68  */
  assign n9930_o = exec[29];
  /* TG68K_ALU.vhd:311:82  */
  assign n9931_o = ~n9930_o;
  /* TG68K_ALU.vhd:311:60  */
  assign n9932_o = n9931_o & n9929_o;
  /* TG68K_ALU.vhd:312:38  */
  assign n9933_o = ~long_start;
  /* TG68K_ALU.vhd:312:59  */
  assign n9935_o = exe_datatype == 2'b00;
  /* TG68K_ALU.vhd:312:43  */
  assign n9936_o = n9935_o & n9933_o;
  /* TG68K_ALU.vhd:312:73  */
  assign n9937_o = exec[50];
  /* TG68K_ALU.vhd:312:81  */
  assign n9938_o = ~n9937_o;
  /* TG68K_ALU.vhd:312:65  */
  assign n9939_o = n9938_o & n9936_o;
  /* TG68K_ALU.vhd:314:41  */
  assign n9940_o = ~long_start;
  /* TG68K_ALU.vhd:314:62  */
  assign n9942_o = exe_datatype == 2'b10;
  /* TG68K_ALU.vhd:314:46  */
  assign n9943_o = n9942_o & n9940_o;
  /* TG68K_ALU.vhd:314:77  */
  assign n9944_o = exec[47];
  /* TG68K_ALU.vhd:314:93  */
  assign n9945_o = exec[46];
  /* TG68K_ALU.vhd:314:86  */
  assign n9946_o = n9944_o | n9945_o;
  /* TG68K_ALU.vhd:314:103  */
  assign n9947_o = n9946_o | movem_presub;
  /* TG68K_ALU.vhd:314:68  */
  assign n9948_o = n9947_o & n9943_o;
  /* TG68K_ALU.vhd:315:40  */
  assign n9949_o = exec[69];
  /* TG68K_ALU.vhd:315:33  */
  assign n9952_o = n9949_o ? 32'b00000000000000000000000000000110 : 32'b00000000000000000000000000000100;
  /* TG68K_ALU.vhd:314:25  */
  assign n9954_o = n9948_o ? n9952_o : 32'b00000000000000000000000000000010;
  /* TG68K_ALU.vhd:312:25  */
  assign n9956_o = n9939_o ? 32'b00000000000000000000000000000001 : n9954_o;
  /* TG68K_ALU.vhd:324:33  */
  assign n9957_o = exec[28];
  /* TG68K_ALU.vhd:324:59  */
  assign n9958_o = n12821_q[4];
  /* TG68K_ALU.vhd:324:50  */
  assign n9959_o = n9958_o & n9957_o;
  /* TG68K_ALU.vhd:324:75  */
  assign n9960_o = exec[31];
  /* TG68K_ALU.vhd:324:68  */
  assign n9961_o = n9959_o | n9960_o;
  /* TG68K_ALU.vhd:324:25  */
  assign n9963_o = n9961_o ? 1'b1 : 1'b0;
  /* TG68K_ALU.vhd:327:41  */
  assign n9964_o = exec[56];
  /* TG68K_ALU.vhd:311:17  */
  assign n9965_o = n9932_o ? n9956_o : op2out;
  /* TG68K_ALU.vhd:311:17  */
  assign n9966_o = n9932_o ? n9916_o : n9964_o;
  /* TG68K_ALU.vhd:311:17  */
  assign n9967_o = n9932_o ? 1'b0 : n9963_o;
  /* TG68KdotC_Kernel.vhd:1407:33  */
  assign n9968_o = n9965_o[15:0];
  /* TG68K_ALU.vhd:309:17  */
  assign n9969_o = n9918_o ? n9925_o : n9968_o;
  assign n9970_o = n9965_o[31:16];
  /* TG68KdotC_Kernel.vhd:1407:33  */
  assign n9971_o = op2out[31:16];
  /* TG68K_ALU.vhd:309:17  */
  assign n9972_o = n9918_o ? n9971_o : n9970_o;
  /* TG68K_ALU.vhd:309:17  */
  assign n9974_o = n9918_o ? n9916_o : n9966_o;
  /* TG68K_ALU.vhd:309:17  */
  assign n9975_o = n9918_o ? 1'b0 : n9967_o;
  /* TG68K_ALU.vhd:331:24  */
  assign n9976_o = exec[69];
  /* TG68K_ALU.vhd:331:43  */
  assign n9977_o = n9976_o | check_aligned;
  /* TG68K_ALU.vhd:332:36  */
  assign n9978_o = ~movem_presub;
  /* TG68K_ALU.vhd:333:64  */
  assign n9979_o = ~long_start;
  /* TG68K_ALU.vhd:333:48  */
  assign n9980_o = n9979_o & non_aligned;
  /* TG68KdotC_Kernel.vhd:1289:1  */
  assign n9982_o = {n9972_o, n9969_o};
  /* TG68K_ALU.vhd:333:25  */
  assign n9983_o = n9980_o ? 32'b00000000000000000000000000000000 : n9982_o;
  /* TG68K_ALU.vhd:337:64  */
  assign n9984_o = ~long_start;
  /* TG68K_ALU.vhd:337:48  */
  assign n9985_o = n9984_o & non_aligned;
  /* TG68K_ALU.vhd:338:44  */
  assign n9987_o = exe_datatype == 2'b10;
  /* TG68K_ALU.vhd:338:27  */
  assign n9990_o = n9987_o ? 32'b00000000000000000000000000001000 : 32'b00000000000000000000000000000100;
  assign n9991_o = {n9972_o, n9969_o};
  /* TG68K_ALU.vhd:337:25  */
  assign n9992_o = n9985_o ? n9990_o : n9991_o;
  /* TG68K_ALU.vhd:332:19  */
  assign n9993_o = n9978_o ? n9983_o : n9992_o;
  assign n9994_o = {n9972_o, n9969_o};
  /* TG68K_ALU.vhd:331:17  */
  assign n9995_o = n9977_o ? n9993_o : n9994_o;
  /* TG68K_ALU.vhd:347:28  */
  assign n9996_o = ~opaddsub;
  /* TG68K_ALU.vhd:347:33  */
  assign n9997_o = n9996_o | long_start;
  /* TG68K_ALU.vhd:348:43  */
  assign n9999_o = {1'b0, addsub_b};
  /* TG68K_ALU.vhd:348:57  */
  assign n10000_o = c_in[0];
  /* TG68K_ALU.vhd:348:52  */
  assign n10001_o = {n9999_o, n10000_o};
  /* TG68K_ALU.vhd:350:48  */
  assign n10003_o = {1'b0, addsub_b};
  /* TG68K_ALU.vhd:350:62  */
  assign n10004_o = c_in[0];
  /* TG68K_ALU.vhd:350:57  */
  assign n10005_o = {n10003_o, n10004_o};
  /* TG68K_ALU.vhd:350:40  */
  assign n10006_o = ~n10005_o;
  /* TG68K_ALU.vhd:347:17  */
  assign n10007_o = n9997_o ? n10001_o : n10006_o;
  /* TG68K_ALU.vhd:352:36  */
  assign n10009_o = {1'b0, addsub_a};
  /* TG68K_ALU.vhd:352:57  */
  assign n10010_o = notaddsub_b[0];
  /* TG68K_ALU.vhd:352:45  */
  assign n10011_o = {n10009_o, n10010_o};
  /* TG68K_ALU.vhd:352:61  */
  assign n10012_o = n10011_o + notaddsub_b;
  /* TG68K_ALU.vhd:353:38  */
  assign n10013_o = add_result[9];
  /* TG68K_ALU.vhd:353:54  */
  assign n10014_o = addsub_a[8];
  /* TG68K_ALU.vhd:353:42  */
  assign n10015_o = n10013_o ^ n10014_o;
  /* TG68K_ALU.vhd:353:70  */
  assign n10016_o = addsub_b[8];
  /* TG68K_ALU.vhd:353:58  */
  assign n10017_o = n10015_o ^ n10016_o;
  /* TG68K_ALU.vhd:354:38  */
  assign n10018_o = add_result[17];
  /* TG68K_ALU.vhd:354:55  */
  assign n10019_o = addsub_a[16];
  /* TG68K_ALU.vhd:354:43  */
  assign n10020_o = n10018_o ^ n10019_o;
  /* TG68K_ALU.vhd:354:72  */
  assign n10021_o = addsub_b[16];
  /* TG68K_ALU.vhd:354:60  */
  assign n10022_o = n10020_o ^ n10021_o;
  /* TG68K_ALU.vhd:355:38  */
  assign n10023_o = add_result[33];
  /* TG68K_ALU.vhd:356:39  */
  assign n10024_o = add_result[32:1];
  /* TG68K_ALU.vhd:357:39  */
  assign n10025_o = c_in[1];
  /* TG68K_ALU.vhd:357:57  */
  assign n10026_o = add_result[8];
  /* TG68K_ALU.vhd:357:43  */
  assign n10027_o = n10025_o ^ n10026_o;
  /* TG68K_ALU.vhd:357:73  */
  assign n10028_o = addsub_a[7];
  /* TG68K_ALU.vhd:357:61  */
  assign n10029_o = n10027_o ^ n10028_o;
  /* TG68K_ALU.vhd:357:89  */
  assign n10030_o = addsub_b[7];
  /* TG68K_ALU.vhd:357:77  */
  assign n10031_o = n10029_o ^ n10030_o;
  /* TG68K_ALU.vhd:358:39  */
  assign n10032_o = c_in[2];
  /* TG68K_ALU.vhd:358:57  */
  assign n10033_o = add_result[16];
  /* TG68K_ALU.vhd:358:43  */
  assign n10034_o = n10032_o ^ n10033_o;
  /* TG68K_ALU.vhd:358:74  */
  assign n10035_o = addsub_a[15];
  /* TG68K_ALU.vhd:358:62  */
  assign n10036_o = n10034_o ^ n10035_o;
  /* TG68K_ALU.vhd:358:91  */
  assign n10037_o = addsub_b[15];
  /* TG68K_ALU.vhd:358:79  */
  assign n10038_o = n10036_o ^ n10037_o;
  /* TG68K_ALU.vhd:359:39  */
  assign n10039_o = c_in[3];
  /* TG68K_ALU.vhd:359:57  */
  assign n10040_o = add_result[32];
  /* TG68K_ALU.vhd:359:43  */
  assign n10041_o = n10039_o ^ n10040_o;
  /* TG68K_ALU.vhd:359:74  */
  assign n10042_o = addsub_a[31];
  /* TG68K_ALU.vhd:359:62  */
  assign n10043_o = n10041_o ^ n10042_o;
  /* TG68K_ALU.vhd:359:91  */
  assign n10044_o = addsub_b[31];
  /* TG68K_ALU.vhd:359:79  */
  assign n10045_o = n10043_o ^ n10044_o;
  /* TG68K_ALU.vhd:360:30  */
  assign n10046_o = c_in[3:1];
  /* TG68K_ALU.vhd:370:32  */
  assign n10050_o = c_in[1];
  /* TG68K_ALU.vhd:370:46  */
  assign n10051_o = add_result[8:0];
  /* TG68K_ALU.vhd:370:35  */
  assign n10052_o = {n10050_o, n10051_o};
  /* TG68K_ALU.vhd:372:38  */
  assign n10053_o = op1out[4];
  /* TG68K_ALU.vhd:372:52  */
  assign n10054_o = op2out[4];
  /* TG68K_ALU.vhd:372:42  */
  assign n10055_o = n10053_o ^ n10054_o;
  /* TG68K_ALU.vhd:372:67  */
  assign n10056_o = bcd_pur[5];
  /* TG68K_ALU.vhd:372:56  */
  assign n10057_o = n10055_o ^ n10056_o;
  /* TG68K_ALU.vhd:373:17  */
  assign n10060_o = halve_carry ? 4'b0110 : 4'b0000;
  /* TG68K_ALU.vhd:376:27  */
  assign n10063_o = bcd_pur[9];
  /* TG68KdotC_Kernel.vhd:217:16  */
  assign n10065_o = n10061_o[7:4];
  /* TG68K_ALU.vhd:376:17  */
  assign n10066_o = n10063_o ? 4'b0110 : n10065_o;
  /* TG68KdotC_Kernel.vhd:174:16  */
  assign n10067_o = n10061_o[8];
  /* TG68K_ALU.vhd:379:24  */
  assign n10068_o = exec[12];
  /* TG68K_ALU.vhd:380:47  */
  assign n10069_o = bcd_pur[8];
  /* TG68K_ALU.vhd:380:36  */
  assign n10070_o = ~n10069_o;
  /* TG68K_ALU.vhd:380:60  */
  assign n10071_o = bcd_a[7];
  /* TG68K_ALU.vhd:380:51  */
  assign n10072_o = n10070_o & n10071_o;
  /* TG68K_ALU.vhd:382:41  */
  assign n10073_o = bcd_pur[9:1];
  /* TG68K_ALU.vhd:382:54  */
  assign n10074_o = n10073_o + bcd_kor;
  /* TG68K_ALU.vhd:383:36  */
  assign n10075_o = bcd_pur[4];
  /* TG68K_ALU.vhd:383:52  */
  assign n10076_o = bcd_pur[3];
  /* TG68K_ALU.vhd:383:66  */
  assign n10077_o = bcd_pur[2];
  /* TG68K_ALU.vhd:383:56  */
  assign n10078_o = n10076_o | n10077_o;
  /* TG68K_ALU.vhd:383:40  */
  assign n10079_o = n10075_o & n10078_o;
  /* TG68K_ALU.vhd:383:25  */
  assign n10081_o = n10079_o ? 4'b0110 : n10060_o;
  /* TG68K_ALU.vhd:386:36  */
  assign n10082_o = bcd_pur[8];
  /* TG68K_ALU.vhd:386:52  */
  assign n10083_o = bcd_pur[7];
  /* TG68K_ALU.vhd:386:66  */
  assign n10084_o = bcd_pur[6];
  /* TG68K_ALU.vhd:386:56  */
  assign n10085_o = n10083_o | n10084_o;
  /* TG68K_ALU.vhd:386:81  */
  assign n10086_o = bcd_pur[5];
  /* TG68K_ALU.vhd:386:96  */
  assign n10087_o = bcd_pur[4];
  /* TG68K_ALU.vhd:386:85  */
  assign n10088_o = n10086_o & n10087_o;
  /* TG68K_ALU.vhd:386:112  */
  assign n10089_o = bcd_pur[3];
  /* TG68K_ALU.vhd:386:126  */
  assign n10090_o = bcd_pur[2];
  /* TG68K_ALU.vhd:386:116  */
  assign n10091_o = n10089_o | n10090_o;
  /* TG68K_ALU.vhd:386:100  */
  assign n10092_o = n10088_o & n10091_o;
  /* TG68K_ALU.vhd:386:70  */
  assign n10093_o = n10085_o | n10092_o;
  /* TG68K_ALU.vhd:386:40  */
  assign n10094_o = n10082_o & n10093_o;
  /* TG68K_ALU.vhd:386:25  */
  assign n10096_o = n10094_o ? 4'b0110 : n10066_o;
  /* TG68K_ALU.vhd:390:43  */
  assign n10097_o = bcd_pur[8];
  /* TG68K_ALU.vhd:390:60  */
  assign n10098_o = bcd_a[7];
  /* TG68K_ALU.vhd:390:51  */
  assign n10099_o = ~n10098_o;
  /* TG68K_ALU.vhd:390:47  */
  assign n10100_o = n10097_o & n10099_o;
  /* TG68K_ALU.vhd:392:41  */
  assign n10101_o = bcd_pur[9:1];
  /* TG68K_ALU.vhd:392:54  */
  assign n10102_o = n10101_o - bcd_kor;
  assign n10103_o = {n10096_o, n10081_o};
  assign n10104_o = {n10066_o, n10060_o};
  /* TG68K_ALU.vhd:379:17  */
  assign n10105_o = n10068_o ? n10103_o : n10104_o;
  /* TG68K_ALU.vhd:379:17  */
  assign n10106_o = n10068_o ? n10072_o : n10100_o;
  /* TG68K_ALU.vhd:379:17  */
  assign n10107_o = n10068_o ? n10074_o : n10102_o;
  /* TG68K_ALU.vhd:394:23  */
  assign n10108_o = cpu[1];
  /* TG68K_ALU.vhd:394:17  */
  assign n10110_o = n10108_o ? 1'b0 : n10106_o;
  /* TG68K_ALU.vhd:397:39  */
  assign n10111_o = bcd_pur[9];
  /* TG68K_ALU.vhd:397:51  */
  assign n10112_o = bcd_a[8];
  /* TG68K_ALU.vhd:397:43  */
  assign n10113_o = n10111_o | n10112_o;
  /* TG68K_ALU.vhd:409:44  */
  assign n10118_o = opcode[7:6];
  /* TG68K_ALU.vhd:410:41  */
  assign n10120_o = n10118_o == 2'b01;
  /* TG68K_ALU.vhd:412:41  */
  assign n10122_o = n10118_o == 2'b11;
  assign n10123_o = {n10122_o, n10120_o};
  /* TG68K_ALU.vhd:409:33  */
  always @*
    case (n10123_o)
      2'b10: n10126_o = 1'b0;
      2'b01: n10126_o = 1'b1;
      default: n10126_o = 1'b0;
    endcase
  /* TG68K_ALU.vhd:409:33  */
  always @*
    case (n10123_o)
      2'b10: n10130_o = 1'b1;
      2'b01: n10130_o = 1'b0;
      default: n10130_o = 1'b0;
    endcase
  /* TG68K_ALU.vhd:419:30  */
  assign n10136_o = exe_opcode[8];
  /* TG68K_ALU.vhd:419:33  */
  assign n10137_o = ~n10136_o;
  /* TG68K_ALU.vhd:420:38  */
  assign n10138_o = exe_opcode[5:4];
  /* TG68K_ALU.vhd:420:50  */
  assign n10140_o = n10138_o == 2'b00;
  /* TG68K_ALU.vhd:421:53  */
  assign n10141_o = sndopc[4:0];
  /* TG68K_ALU.vhd:423:58  */
  assign n10142_o = sndopc[2:0];
  /* TG68K_ALU.vhd:423:51  */
  assign n10144_o = {2'b00, n10142_o};
  /* TG68K_ALU.vhd:420:25  */
  assign n10145_o = n10140_o ? n10141_o : n10144_o;
  /* TG68K_ALU.vhd:426:38  */
  assign n10146_o = exe_opcode[5:4];
  /* TG68K_ALU.vhd:426:50  */
  assign n10148_o = n10146_o == 2'b00;
  /* TG68K_ALU.vhd:427:53  */
  assign n10149_o = reg_qb[4:0];
  /* TG68K_ALU.vhd:429:58  */
  assign n10150_o = reg_qb[2:0];
  /* TG68K_ALU.vhd:429:51  */
  assign n10152_o = {2'b00, n10150_o};
  /* TG68K_ALU.vhd:426:25  */
  assign n10153_o = n10148_o ? n10149_o : n10152_o;
  /* TG68K_ALU.vhd:419:17  */
  assign n10154_o = n10137_o ? n10145_o : n10153_o;
  /* TG68K_ALU.vhd:435:65  */
  assign n10160_o = ~one_bit_in;
  /* TG68K_ALU.vhd:435:61  */
  assign n10161_o = bchg & n10160_o;
  /* TG68K_ALU.vhd:435:81  */
  assign n10162_o = n10161_o | bset;
  /* TG68K_ALU.vhd:456:42  */
  assign n10168_o = opcode[5:4];
  /* TG68K_ALU.vhd:456:55  */
  assign n10170_o = n10168_o == 2'b00;
  /* TG68K_ALU.vhd:456:33  */
  assign n10173_o = n10170_o ? 1'b1 : 1'b0;
  /* TG68K_ALU.vhd:459:44  */
  assign n10175_o = opcode[10:8];
  /* TG68K_ALU.vhd:460:41  */
  assign n10177_o = n10175_o == 3'b010;
  /* TG68K_ALU.vhd:461:41  */
  assign n10179_o = n10175_o == 3'b011;
  /* TG68K_ALU.vhd:463:41  */
  assign n10181_o = n10175_o == 3'b101;
  /* TG68K_ALU.vhd:464:41  */
  assign n10183_o = n10175_o == 3'b110;
  /* TG68K_ALU.vhd:465:41  */
  assign n10185_o = n10175_o == 3'b111;
  assign n10186_o = {n10185_o, n10183_o, n10181_o, n10179_o, n10177_o};
  /* TG68K_ALU.vhd:459:33  */
  always @*
    case (n10186_o)
      5'b10000: n10189_o = 1'b0;
      5'b01000: n10189_o = 1'b1;
      5'b00100: n10189_o = 1'b0;
      5'b00010: n10189_o = 1'b0;
      5'b00001: n10189_o = 1'b0;
      default: n10189_o = 1'b0;
    endcase
  /* TG68K_ALU.vhd:459:33  */
  always @*
    case (n10186_o)
      5'b10000: n10193_o = 1'b0;
      5'b01000: n10193_o = 1'b0;
      5'b00100: n10193_o = 1'b0;
      5'b00010: n10193_o = 1'b0;
      5'b00001: n10193_o = 1'b1;
      default: n10193_o = 1'b0;
    endcase
  /* TG68K_ALU.vhd:459:33  */
  always @*
    case (n10186_o)
      5'b10000: n10197_o = 1'b1;
      5'b01000: n10197_o = 1'b0;
      5'b00100: n10197_o = 1'b0;
      5'b00010: n10197_o = 1'b0;
      5'b00001: n10197_o = 1'b0;
      default: n10197_o = 1'b0;
    endcase
  /* TG68K_ALU.vhd:459:33  */
  always @*
    case (n10186_o)
      5'b10000: n10201_o = 1'b0;
      5'b01000: n10201_o = 1'b0;
      5'b00100: n10201_o = 1'b0;
      5'b00010: n10201_o = 1'b1;
      5'b00001: n10201_o = 1'b0;
      default: n10201_o = 1'b0;
    endcase
  /* TG68K_ALU.vhd:459:33  */
  always @*
    case (n10186_o)
      5'b10000: n10205_o = 1'b0;
      5'b01000: n10205_o = 1'b0;
      5'b00100: n10205_o = 1'b1;
      5'b00010: n10205_o = 1'b0;
      5'b00001: n10205_o = 1'b0;
      default: n10205_o = 1'b0;
    endcase
  /* TG68K_ALU.vhd:459:33  */
  always @*
    case (n10186_o)
      5'b10000: n10208_o = 1'b1;
      5'b01000: n10208_o = n10173_o;
      5'b00100: n10208_o = n10173_o;
      5'b00010: n10208_o = n10173_o;
      5'b00001: n10208_o = n10173_o;
      default: n10208_o = n10173_o;
    endcase
  /* TG68K_ALU.vhd:469:42  */
  assign n10209_o = opcode[4:3];
  /* TG68K_ALU.vhd:469:54  */
  assign n10211_o = n10209_o == 2'b00;
  /* TG68K_ALU.vhd:469:33  */
  assign n10214_o = n10211_o ? 1'b1 : 1'b0;
  /* TG68K_ALU.vhd:472:53  */
  assign n10216_o = result[39:32];
  /* TG68K_ALU.vhd:490:38  */
  assign n10234_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10236_o = $unsigned(5'b00000) > $unsigned(n10234_o);
  assign n10239_o = reg_qb[0];
  assign n10240_o = bf_set2[0];
  /* TG68K_ALU.vhd:476:17  */
  assign n10241_o = bf_ins ? n10239_o : n10240_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10242_o = n10236_o ? 1'b0 : n10241_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10247_o = n10236_o ? 1'b1 : 1'b0;
  /* TG68K_ALU.vhd:490:38  */
  assign n10250_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10252_o = $unsigned(5'b00001) > $unsigned(n10250_o);
  assign n10255_o = reg_qb[1];
  assign n10256_o = bf_set2[1];
  /* TG68K_ALU.vhd:476:17  */
  assign n10257_o = bf_ins ? n10255_o : n10256_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10258_o = n10252_o ? 1'b0 : n10257_o;
  assign n10262_o = n10248_o[1];
  /* TG68K_ALU.vhd:490:25  */
  assign n10263_o = n10252_o ? 1'b1 : n10262_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10265_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10267_o = $unsigned(5'b00010) > $unsigned(n10265_o);
  assign n10270_o = reg_qb[2];
  assign n10271_o = bf_set2[2];
  /* TG68K_ALU.vhd:476:17  */
  assign n10272_o = bf_ins ? n10270_o : n10271_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10273_o = n10267_o ? 1'b0 : n10272_o;
  assign n10277_o = n10248_o[2];
  /* TG68K_ALU.vhd:490:25  */
  assign n10278_o = n10267_o ? 1'b1 : n10277_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10280_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10282_o = $unsigned(5'b00011) > $unsigned(n10280_o);
  assign n10285_o = reg_qb[3];
  assign n10286_o = bf_set2[3];
  /* TG68K_ALU.vhd:476:17  */
  assign n10287_o = bf_ins ? n10285_o : n10286_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10288_o = n10282_o ? 1'b0 : n10287_o;
  assign n10292_o = n10248_o[3];
  /* TG68K_ALU.vhd:490:25  */
  assign n10293_o = n10282_o ? 1'b1 : n10292_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10295_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10297_o = $unsigned(5'b00100) > $unsigned(n10295_o);
  assign n10300_o = reg_qb[4];
  assign n10301_o = bf_set2[4];
  /* TG68K_ALU.vhd:476:17  */
  assign n10302_o = bf_ins ? n10300_o : n10301_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10303_o = n10297_o ? 1'b0 : n10302_o;
  assign n10307_o = n10248_o[4];
  /* TG68K_ALU.vhd:490:25  */
  assign n10308_o = n10297_o ? 1'b1 : n10307_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10310_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10312_o = $unsigned(5'b00101) > $unsigned(n10310_o);
  assign n10315_o = reg_qb[5];
  assign n10316_o = bf_set2[5];
  /* TG68K_ALU.vhd:476:17  */
  assign n10317_o = bf_ins ? n10315_o : n10316_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10318_o = n10312_o ? 1'b0 : n10317_o;
  assign n10322_o = n10248_o[5];
  /* TG68K_ALU.vhd:490:25  */
  assign n10323_o = n10312_o ? 1'b1 : n10322_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10325_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10327_o = $unsigned(5'b00110) > $unsigned(n10325_o);
  assign n10330_o = reg_qb[6];
  assign n10331_o = bf_set2[6];
  /* TG68K_ALU.vhd:476:17  */
  assign n10332_o = bf_ins ? n10330_o : n10331_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10333_o = n10327_o ? 1'b0 : n10332_o;
  assign n10337_o = n10248_o[6];
  /* TG68K_ALU.vhd:490:25  */
  assign n10338_o = n10327_o ? 1'b1 : n10337_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10340_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10342_o = $unsigned(5'b00111) > $unsigned(n10340_o);
  assign n10345_o = reg_qb[7];
  assign n10346_o = bf_set2[7];
  /* TG68K_ALU.vhd:476:17  */
  assign n10347_o = bf_ins ? n10345_o : n10346_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10348_o = n10342_o ? 1'b0 : n10347_o;
  assign n10352_o = n10248_o[7];
  /* TG68K_ALU.vhd:490:25  */
  assign n10353_o = n10342_o ? 1'b1 : n10352_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10355_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10357_o = $unsigned(5'b01000) > $unsigned(n10355_o);
  assign n10360_o = reg_qb[8];
  assign n10361_o = bf_set2[8];
  /* TG68K_ALU.vhd:476:17  */
  assign n10362_o = bf_ins ? n10360_o : n10361_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10363_o = n10357_o ? 1'b0 : n10362_o;
  assign n10367_o = n10248_o[8];
  /* TG68K_ALU.vhd:490:25  */
  assign n10368_o = n10357_o ? 1'b1 : n10367_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10370_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10372_o = $unsigned(5'b01001) > $unsigned(n10370_o);
  assign n10375_o = reg_qb[9];
  assign n10376_o = bf_set2[9];
  /* TG68K_ALU.vhd:476:17  */
  assign n10377_o = bf_ins ? n10375_o : n10376_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10378_o = n10372_o ? 1'b0 : n10377_o;
  assign n10382_o = n10248_o[9];
  /* TG68K_ALU.vhd:490:25  */
  assign n10383_o = n10372_o ? 1'b1 : n10382_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10385_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10387_o = $unsigned(5'b01010) > $unsigned(n10385_o);
  assign n10390_o = reg_qb[10];
  assign n10391_o = bf_set2[10];
  /* TG68K_ALU.vhd:476:17  */
  assign n10392_o = bf_ins ? n10390_o : n10391_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10393_o = n10387_o ? 1'b0 : n10392_o;
  assign n10397_o = n10248_o[10];
  /* TG68K_ALU.vhd:490:25  */
  assign n10398_o = n10387_o ? 1'b1 : n10397_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10400_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10402_o = $unsigned(5'b01011) > $unsigned(n10400_o);
  assign n10405_o = reg_qb[11];
  assign n10406_o = bf_set2[11];
  /* TG68K_ALU.vhd:476:17  */
  assign n10407_o = bf_ins ? n10405_o : n10406_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10408_o = n10402_o ? 1'b0 : n10407_o;
  assign n10412_o = n10248_o[11];
  /* TG68K_ALU.vhd:490:25  */
  assign n10413_o = n10402_o ? 1'b1 : n10412_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10415_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10417_o = $unsigned(5'b01100) > $unsigned(n10415_o);
  assign n10420_o = reg_qb[12];
  assign n10421_o = bf_set2[12];
  /* TG68K_ALU.vhd:476:17  */
  assign n10422_o = bf_ins ? n10420_o : n10421_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10423_o = n10417_o ? 1'b0 : n10422_o;
  assign n10427_o = n10248_o[12];
  /* TG68K_ALU.vhd:490:25  */
  assign n10428_o = n10417_o ? 1'b1 : n10427_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10430_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10432_o = $unsigned(5'b01101) > $unsigned(n10430_o);
  assign n10435_o = reg_qb[13];
  assign n10436_o = bf_set2[13];
  /* TG68K_ALU.vhd:476:17  */
  assign n10437_o = bf_ins ? n10435_o : n10436_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10438_o = n10432_o ? 1'b0 : n10437_o;
  assign n10442_o = n10248_o[13];
  /* TG68K_ALU.vhd:490:25  */
  assign n10443_o = n10432_o ? 1'b1 : n10442_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10445_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10447_o = $unsigned(5'b01110) > $unsigned(n10445_o);
  assign n10450_o = reg_qb[14];
  assign n10451_o = bf_set2[14];
  /* TG68K_ALU.vhd:476:17  */
  assign n10452_o = bf_ins ? n10450_o : n10451_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10453_o = n10447_o ? 1'b0 : n10452_o;
  assign n10457_o = n10248_o[14];
  /* TG68K_ALU.vhd:490:25  */
  assign n10458_o = n10447_o ? 1'b1 : n10457_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10460_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10462_o = $unsigned(5'b01111) > $unsigned(n10460_o);
  assign n10465_o = reg_qb[15];
  assign n10466_o = bf_set2[15];
  /* TG68K_ALU.vhd:476:17  */
  assign n10467_o = bf_ins ? n10465_o : n10466_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10468_o = n10462_o ? 1'b0 : n10467_o;
  assign n10472_o = n10248_o[15];
  /* TG68K_ALU.vhd:490:25  */
  assign n10473_o = n10462_o ? 1'b1 : n10472_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10475_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10477_o = $unsigned(5'b10000) > $unsigned(n10475_o);
  assign n10480_o = reg_qb[16];
  assign n10481_o = bf_set2[16];
  /* TG68K_ALU.vhd:476:17  */
  assign n10482_o = bf_ins ? n10480_o : n10481_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10483_o = n10477_o ? 1'b0 : n10482_o;
  assign n10487_o = n10248_o[16];
  /* TG68K_ALU.vhd:490:25  */
  assign n10488_o = n10477_o ? 1'b1 : n10487_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10490_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10492_o = $unsigned(5'b10001) > $unsigned(n10490_o);
  assign n10495_o = reg_qb[17];
  assign n10496_o = bf_set2[17];
  /* TG68K_ALU.vhd:476:17  */
  assign n10497_o = bf_ins ? n10495_o : n10496_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10498_o = n10492_o ? 1'b0 : n10497_o;
  assign n10502_o = n10248_o[17];
  /* TG68K_ALU.vhd:490:25  */
  assign n10503_o = n10492_o ? 1'b1 : n10502_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10505_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10507_o = $unsigned(5'b10010) > $unsigned(n10505_o);
  assign n10510_o = reg_qb[18];
  assign n10511_o = bf_set2[18];
  /* TG68K_ALU.vhd:476:17  */
  assign n10512_o = bf_ins ? n10510_o : n10511_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10513_o = n10507_o ? 1'b0 : n10512_o;
  assign n10517_o = n10248_o[18];
  /* TG68K_ALU.vhd:490:25  */
  assign n10518_o = n10507_o ? 1'b1 : n10517_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10520_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10522_o = $unsigned(5'b10011) > $unsigned(n10520_o);
  assign n10525_o = reg_qb[19];
  assign n10526_o = bf_set2[19];
  /* TG68K_ALU.vhd:476:17  */
  assign n10527_o = bf_ins ? n10525_o : n10526_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10528_o = n10522_o ? 1'b0 : n10527_o;
  assign n10532_o = n10248_o[19];
  /* TG68K_ALU.vhd:490:25  */
  assign n10533_o = n10522_o ? 1'b1 : n10532_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10535_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10537_o = $unsigned(5'b10100) > $unsigned(n10535_o);
  assign n10540_o = reg_qb[20];
  assign n10541_o = bf_set2[20];
  /* TG68K_ALU.vhd:476:17  */
  assign n10542_o = bf_ins ? n10540_o : n10541_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10543_o = n10537_o ? 1'b0 : n10542_o;
  assign n10547_o = n10248_o[20];
  /* TG68K_ALU.vhd:490:25  */
  assign n10548_o = n10537_o ? 1'b1 : n10547_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10550_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10552_o = $unsigned(5'b10101) > $unsigned(n10550_o);
  assign n10555_o = reg_qb[21];
  assign n10556_o = bf_set2[21];
  /* TG68K_ALU.vhd:476:17  */
  assign n10557_o = bf_ins ? n10555_o : n10556_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10558_o = n10552_o ? 1'b0 : n10557_o;
  assign n10562_o = n10248_o[21];
  /* TG68K_ALU.vhd:490:25  */
  assign n10563_o = n10552_o ? 1'b1 : n10562_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10565_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10567_o = $unsigned(5'b10110) > $unsigned(n10565_o);
  assign n10570_o = reg_qb[22];
  assign n10571_o = bf_set2[22];
  /* TG68K_ALU.vhd:476:17  */
  assign n10572_o = bf_ins ? n10570_o : n10571_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10573_o = n10567_o ? 1'b0 : n10572_o;
  assign n10577_o = n10248_o[22];
  /* TG68K_ALU.vhd:490:25  */
  assign n10578_o = n10567_o ? 1'b1 : n10577_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10580_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10582_o = $unsigned(5'b10111) > $unsigned(n10580_o);
  assign n10585_o = reg_qb[23];
  assign n10586_o = bf_set2[23];
  /* TG68K_ALU.vhd:476:17  */
  assign n10587_o = bf_ins ? n10585_o : n10586_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10588_o = n10582_o ? 1'b0 : n10587_o;
  assign n10592_o = n10248_o[23];
  /* TG68K_ALU.vhd:490:25  */
  assign n10593_o = n10582_o ? 1'b1 : n10592_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10595_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10597_o = $unsigned(5'b11000) > $unsigned(n10595_o);
  assign n10600_o = reg_qb[24];
  assign n10601_o = bf_set2[24];
  /* TG68K_ALU.vhd:476:17  */
  assign n10602_o = bf_ins ? n10600_o : n10601_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10603_o = n10597_o ? 1'b0 : n10602_o;
  assign n10607_o = n10248_o[24];
  /* TG68K_ALU.vhd:490:25  */
  assign n10608_o = n10597_o ? 1'b1 : n10607_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10610_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10612_o = $unsigned(5'b11001) > $unsigned(n10610_o);
  assign n10615_o = reg_qb[25];
  assign n10616_o = bf_set2[25];
  /* TG68K_ALU.vhd:476:17  */
  assign n10617_o = bf_ins ? n10615_o : n10616_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10618_o = n10612_o ? 1'b0 : n10617_o;
  assign n10622_o = n10248_o[25];
  /* TG68K_ALU.vhd:490:25  */
  assign n10623_o = n10612_o ? 1'b1 : n10622_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10625_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10627_o = $unsigned(5'b11010) > $unsigned(n10625_o);
  assign n10630_o = reg_qb[26];
  assign n10631_o = bf_set2[26];
  /* TG68K_ALU.vhd:476:17  */
  assign n10632_o = bf_ins ? n10630_o : n10631_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10633_o = n10627_o ? 1'b0 : n10632_o;
  assign n10637_o = n10248_o[26];
  /* TG68K_ALU.vhd:490:25  */
  assign n10638_o = n10627_o ? 1'b1 : n10637_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10640_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10642_o = $unsigned(5'b11011) > $unsigned(n10640_o);
  assign n10645_o = reg_qb[27];
  assign n10646_o = bf_set2[27];
  /* TG68K_ALU.vhd:476:17  */
  assign n10647_o = bf_ins ? n10645_o : n10646_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10648_o = n10642_o ? 1'b0 : n10647_o;
  assign n10652_o = n10248_o[27];
  /* TG68K_ALU.vhd:490:25  */
  assign n10653_o = n10642_o ? 1'b1 : n10652_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10655_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10657_o = $unsigned(5'b11100) > $unsigned(n10655_o);
  assign n10660_o = reg_qb[28];
  assign n10661_o = bf_set2[28];
  /* TG68K_ALU.vhd:476:17  */
  assign n10662_o = bf_ins ? n10660_o : n10661_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10663_o = n10657_o ? 1'b0 : n10662_o;
  assign n10667_o = n10248_o[28];
  /* TG68K_ALU.vhd:490:25  */
  assign n10668_o = n10657_o ? 1'b1 : n10667_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10670_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10672_o = $unsigned(5'b11101) > $unsigned(n10670_o);
  assign n10675_o = reg_qb[29];
  assign n10676_o = bf_set2[29];
  /* TG68K_ALU.vhd:476:17  */
  assign n10677_o = bf_ins ? n10675_o : n10676_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10678_o = n10672_o ? 1'b0 : n10677_o;
  assign n10682_o = n10248_o[29];
  /* TG68K_ALU.vhd:490:25  */
  assign n10683_o = n10672_o ? 1'b1 : n10682_o;
  /* TG68K_ALU.vhd:490:38  */
  assign n10685_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10687_o = $unsigned(5'b11110) > $unsigned(n10685_o);
  assign n10690_o = reg_qb[30];
  assign n10691_o = bf_set2[30];
  /* TG68K_ALU.vhd:476:17  */
  assign n10692_o = bf_ins ? n10690_o : n10691_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10693_o = n10687_o ? 1'b0 : n10692_o;
  assign n10694_o = reg_qb[31];
  assign n10695_o = bf_set2[31];
  /* TG68K_ALU.vhd:476:17  */
  assign n10696_o = bf_ins ? n10694_o : n10695_o;
  assign n10697_o = n10248_o[30];
  /* TG68K_ALU.vhd:490:25  */
  assign n10698_o = n10687_o ? 1'b1 : n10697_o;
  assign n10699_o = n10248_o[31];
  /* TG68K_ALU.vhd:490:38  */
  assign n10700_o = bf_width[4:0];
  /* TG68K_ALU.vhd:490:29  */
  assign n10702_o = $unsigned(5'b11111) > $unsigned(n10700_o);
  /* TG68K_ALU.vhd:490:25  */
  assign n10705_o = n10702_o ? 1'b0 : n10696_o;
  /* TG68K_ALU.vhd:490:25  */
  assign n10706_o = n10702_o ? 1'b1 : n10699_o;
  /* TG68K_ALU.vhd:496:37  */
  assign n10708_o = bf_width[4:0];  // trunc
  /* TG68K_ALU.vhd:497:32  */
  assign n10711_o = bf_nflag & bf_exts;
  /* TG68K_ALU.vhd:498:47  */
  assign n10712_o = datareg | unshifted_bitmask;
  /* TG68K_ALU.vhd:497:17  */
  assign n10713_o = n10711_o ? n10712_o : datareg;
  /* TG68K_ALU.vhd:504:30  */
  assign n10714_o = bf_loffset[4];
  /* TG68K_ALU.vhd:505:57  */
  assign n10715_o = unshifted_bitmask[15:0];
  /* TG68K_ALU.vhd:505:88  */
  assign n10716_o = unshifted_bitmask[31:16];
  /* TG68K_ALU.vhd:505:70  */
  assign n10717_o = {n10715_o, n10716_o};
  /* TG68K_ALU.vhd:504:17  */
  assign n10718_o = n10714_o ? n10717_o : unshifted_bitmask;
  /* TG68K_ALU.vhd:509:30  */
  assign n10719_o = bf_loffset[3];
  /* TG68K_ALU.vhd:510:64  */
  assign n10720_o = bitmaskmux3[23:0];
  /* TG68K_ALU.vhd:510:89  */
  assign n10721_o = bitmaskmux3[31:24];
  /* TG68K_ALU.vhd:510:77  */
  assign n10722_o = {n10720_o, n10721_o};
  /* TG68K_ALU.vhd:509:17  */
  assign n10723_o = n10719_o ? n10722_o : bitmaskmux3;
  /* TG68K_ALU.vhd:514:30  */
  assign n10724_o = bf_loffset[2];
  /* TG68K_ALU.vhd:515:51  */
  assign n10726_o = {bitmaskmux2, 4'b1111};
  /* TG68K_ALU.vhd:517:71  */
  assign n10727_o = bitmaskmux2[31:28];
  assign n10728_o = n10726_o[3:0];
  /* TG68K_ALU.vhd:516:25  */
  assign n10729_o = bf_d32 ? n10727_o : n10728_o;
  assign n10730_o = n10726_o[35:4];
  /* TG68K_ALU.vhd:520:46  */
  assign n10732_o = {4'b1111, bitmaskmux2};
  assign n10733_o = {n10730_o, n10729_o};
  /* TG68K_ALU.vhd:514:17  */
  assign n10734_o = n10724_o ? n10733_o : n10732_o;
  /* TG68K_ALU.vhd:522:30  */
  assign n10735_o = bf_loffset[1];
  /* TG68K_ALU.vhd:523:51  */
  assign n10737_o = {bitmaskmux1, 2'b11};
  /* TG68K_ALU.vhd:525:71  */
  assign n10738_o = bitmaskmux1[31:30];
  assign n10739_o = n10737_o[1:0];
  /* TG68K_ALU.vhd:524:25  */
  assign n10740_o = bf_d32 ? n10738_o : n10739_o;
  assign n10741_o = n10737_o[37:2];
  /* TG68K_ALU.vhd:528:44  */
  assign n10743_o = {2'b11, bitmaskmux1};
  assign n10744_o = {n10741_o, n10740_o};
  /* TG68K_ALU.vhd:522:17  */
  assign n10745_o = n10735_o ? n10744_o : n10743_o;
  /* TG68K_ALU.vhd:530:30  */
  assign n10746_o = bf_loffset[0];
  /* TG68K_ALU.vhd:531:47  */
  assign n10748_o = {1'b1, bitmaskmux0};
  /* TG68K_ALU.vhd:531:59  */
  assign n10750_o = {n10748_o, 1'b1};
  /* TG68K_ALU.vhd:533:66  */
  assign n10751_o = bitmaskmux0[31];
  assign n10752_o = n10750_o[0];
  /* TG68K_ALU.vhd:532:25  */
  assign n10753_o = bf_d32 ? n10751_o : n10752_o;
  assign n10754_o = n10750_o[39:1];
  /* TG68K_ALU.vhd:536:48  */
  assign n10756_o = {2'b11, bitmaskmux0};
  assign n10757_o = {n10754_o, n10753_o};
  /* TG68K_ALU.vhd:530:17  */
  assign n10758_o = n10746_o ? n10757_o : n10756_o;
  /* TG68K_ALU.vhd:541:35  */
  assign n10759_o = {bf_ext_in, op2out};
  /* TG68K_ALU.vhd:543:54  */
  assign n10760_o = op2out[7:0];
  assign n10761_o = n10759_o[39:32];
  /* TG68K_ALU.vhd:542:17  */
  assign n10762_o = bf_s32 ? n10760_o : n10761_o;
  assign n10763_o = n10759_o[31:0];
  /* TG68K_ALU.vhd:546:28  */
  assign n10764_o = bf_shift[0];
  /* TG68K_ALU.vhd:547:40  */
  assign n10765_o = shift[0];
  /* TG68K_ALU.vhd:547:49  */
  assign n10766_o = shift[39:1];
  /* TG68K_ALU.vhd:547:43  */
  assign n10767_o = {n10765_o, n10766_o};
  /* TG68K_ALU.vhd:546:17  */
  assign n10768_o = n10764_o ? n10767_o : shift;
  /* TG68K_ALU.vhd:551:28  */
  assign n10769_o = bf_shift[1];
  /* TG68K_ALU.vhd:552:41  */
  assign n10770_o = inmux0[1:0];
  /* TG68K_ALU.vhd:552:60  */
  assign n10771_o = inmux0[39:2];
  /* TG68K_ALU.vhd:552:53  */
  assign n10772_o = {n10770_o, n10771_o};
  /* TG68K_ALU.vhd:551:17  */
  assign n10773_o = n10769_o ? n10772_o : inmux0;
  /* TG68K_ALU.vhd:556:28  */
  assign n10774_o = bf_shift[2];
  /* TG68K_ALU.vhd:557:41  */
  assign n10775_o = inmux1[3:0];
  /* TG68K_ALU.vhd:557:60  */
  assign n10776_o = inmux1[39:4];
  /* TG68K_ALU.vhd:557:53  */
  assign n10777_o = {n10775_o, n10776_o};
  /* TG68K_ALU.vhd:556:17  */
  assign n10778_o = n10774_o ? n10777_o : inmux1;
  /* TG68K_ALU.vhd:561:28  */
  assign n10779_o = bf_shift[3];
  /* TG68K_ALU.vhd:562:41  */
  assign n10780_o = inmux2[7:0];
  /* TG68K_ALU.vhd:562:60  */
  assign n10781_o = inmux2[31:8];
  /* TG68K_ALU.vhd:562:53  */
  assign n10782_o = {n10780_o, n10781_o};
  /* TG68K_ALU.vhd:564:41  */
  assign n10783_o = inmux2[31:0];
  /* TG68K_ALU.vhd:561:17  */
  assign n10784_o = n10779_o ? n10782_o : n10783_o;
  /* TG68K_ALU.vhd:566:28  */
  assign n10785_o = bf_shift[4];
  /* TG68K_ALU.vhd:567:55  */
  assign n10786_o = inmux3[15:0];
  /* TG68K_ALU.vhd:567:75  */
  assign n10787_o = inmux3[31:16];
  /* TG68K_ALU.vhd:567:68  */
  assign n10788_o = {n10786_o, n10787_o};
  /* TG68K_ALU.vhd:566:17  */
  assign n10789_o = n10785_o ? n10788_o : inmux3;
  /* TG68K_ALU.vhd:574:56  */
  assign n10790_o = bf_set2[7:0];
  /* TG68K_ALU.vhd:576:48  */
  assign n10791_o = ~op2out;
  /* TG68K_ALU.vhd:577:49  */
  assign n10792_o = ~bf_ext_in;
  assign n10793_o = {n10792_o, n10791_o};
  assign n10796_o = {n10790_o, bf_set2};
  /* TG68K_ALU.vhd:586:48  */
  assign n10800_o = {bf_ext_in, op1out};
  /* TG68K_ALU.vhd:588:48  */
  assign n10801_o = {bf_ext_in, op2out};
  /* TG68K_ALU.vhd:585:17  */
  assign n10802_o = bf_ins ? n10800_o : n10801_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n10803_o = shifted_bitmask[0];
  /* TG68K_ALU.vhd:592:56  */
  assign n10804_o = result_tmp[0];
  assign n10805_o = n10798_o[0];
  assign n10806_o = n10796_o[0];
  assign n10807_o = n10793_o[0];
  assign n10808_o = n10794_o[0];
  /* TG68K_ALU.vhd:575:17  */
  assign n10809_o = bf_bchg ? n10807_o : n10808_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n10810_o = bf_ins ? n10806_o : n10809_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n10811_o = bf_bset ? n10805_o : n10810_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n10812_o = n10803_o ? n10804_o : n10811_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n10820_o = shifted_bitmask[1];
  /* TG68K_ALU.vhd:592:56  */
  assign n10821_o = result_tmp[1];
  assign n10822_o = n10798_o[1];
  assign n10823_o = n10796_o[1];
  assign n10824_o = n10793_o[1];
  assign n10825_o = n10794_o[1];
  /* TG68K_ALU.vhd:575:17  */
  assign n10826_o = bf_bchg ? n10824_o : n10825_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n10827_o = bf_ins ? n10823_o : n10826_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n10828_o = bf_bset ? n10822_o : n10827_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n10829_o = n10820_o ? n10821_o : n10828_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n10837_o = shifted_bitmask[2];
  /* TG68K_ALU.vhd:592:56  */
  assign n10838_o = result_tmp[2];
  assign n10839_o = n10798_o[2];
  assign n10840_o = n10796_o[2];
  assign n10841_o = n10793_o[2];
  assign n10842_o = n10794_o[2];
  /* TG68K_ALU.vhd:575:17  */
  assign n10843_o = bf_bchg ? n10841_o : n10842_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n10844_o = bf_ins ? n10840_o : n10843_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n10845_o = bf_bset ? n10839_o : n10844_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n10846_o = n10837_o ? n10838_o : n10845_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n10854_o = shifted_bitmask[3];
  /* TG68K_ALU.vhd:592:56  */
  assign n10855_o = result_tmp[3];
  assign n10856_o = n10798_o[3];
  assign n10857_o = n10796_o[3];
  assign n10858_o = n10793_o[3];
  assign n10859_o = n10794_o[3];
  /* TG68K_ALU.vhd:575:17  */
  assign n10860_o = bf_bchg ? n10858_o : n10859_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n10861_o = bf_ins ? n10857_o : n10860_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n10862_o = bf_bset ? n10856_o : n10861_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n10863_o = n10854_o ? n10855_o : n10862_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n10871_o = shifted_bitmask[4];
  /* TG68K_ALU.vhd:592:56  */
  assign n10872_o = result_tmp[4];
  assign n10873_o = n10798_o[4];
  assign n10874_o = n10796_o[4];
  assign n10875_o = n10793_o[4];
  assign n10876_o = n10794_o[4];
  /* TG68K_ALU.vhd:575:17  */
  assign n10877_o = bf_bchg ? n10875_o : n10876_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n10878_o = bf_ins ? n10874_o : n10877_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n10879_o = bf_bset ? n10873_o : n10878_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n10880_o = n10871_o ? n10872_o : n10879_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n10888_o = shifted_bitmask[5];
  /* TG68K_ALU.vhd:592:56  */
  assign n10889_o = result_tmp[5];
  assign n10890_o = n10798_o[5];
  assign n10891_o = n10796_o[5];
  assign n10892_o = n10793_o[5];
  assign n10893_o = n10794_o[5];
  /* TG68K_ALU.vhd:575:17  */
  assign n10894_o = bf_bchg ? n10892_o : n10893_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n10895_o = bf_ins ? n10891_o : n10894_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n10896_o = bf_bset ? n10890_o : n10895_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n10897_o = n10888_o ? n10889_o : n10896_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n10905_o = shifted_bitmask[6];
  /* TG68K_ALU.vhd:592:56  */
  assign n10906_o = result_tmp[6];
  assign n10907_o = n10798_o[6];
  assign n10908_o = n10796_o[6];
  assign n10909_o = n10793_o[6];
  assign n10910_o = n10794_o[6];
  /* TG68K_ALU.vhd:575:17  */
  assign n10911_o = bf_bchg ? n10909_o : n10910_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n10912_o = bf_ins ? n10908_o : n10911_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n10913_o = bf_bset ? n10907_o : n10912_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n10914_o = n10905_o ? n10906_o : n10913_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n10922_o = shifted_bitmask[7];
  /* TG68K_ALU.vhd:592:56  */
  assign n10923_o = result_tmp[7];
  assign n10924_o = n10798_o[7];
  assign n10925_o = n10796_o[7];
  assign n10926_o = n10793_o[7];
  assign n10927_o = n10794_o[7];
  /* TG68K_ALU.vhd:575:17  */
  assign n10928_o = bf_bchg ? n10926_o : n10927_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n10929_o = bf_ins ? n10925_o : n10928_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n10930_o = bf_bset ? n10924_o : n10929_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n10931_o = n10922_o ? n10923_o : n10930_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n10939_o = shifted_bitmask[8];
  /* TG68K_ALU.vhd:592:56  */
  assign n10940_o = result_tmp[8];
  assign n10941_o = n10798_o[8];
  assign n10942_o = n10796_o[8];
  assign n10943_o = n10793_o[8];
  assign n10944_o = n10794_o[8];
  /* TG68K_ALU.vhd:575:17  */
  assign n10945_o = bf_bchg ? n10943_o : n10944_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n10946_o = bf_ins ? n10942_o : n10945_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n10947_o = bf_bset ? n10941_o : n10946_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n10948_o = n10939_o ? n10940_o : n10947_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n10956_o = shifted_bitmask[9];
  /* TG68K_ALU.vhd:592:56  */
  assign n10957_o = result_tmp[9];
  assign n10958_o = n10798_o[9];
  assign n10959_o = n10796_o[9];
  assign n10960_o = n10793_o[9];
  assign n10961_o = n10794_o[9];
  /* TG68K_ALU.vhd:575:17  */
  assign n10962_o = bf_bchg ? n10960_o : n10961_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n10963_o = bf_ins ? n10959_o : n10962_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n10964_o = bf_bset ? n10958_o : n10963_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n10965_o = n10956_o ? n10957_o : n10964_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n10973_o = shifted_bitmask[10];
  /* TG68K_ALU.vhd:592:56  */
  assign n10974_o = result_tmp[10];
  assign n10975_o = n10798_o[10];
  assign n10976_o = n10796_o[10];
  assign n10977_o = n10793_o[10];
  assign n10978_o = n10794_o[10];
  /* TG68K_ALU.vhd:575:17  */
  assign n10979_o = bf_bchg ? n10977_o : n10978_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n10980_o = bf_ins ? n10976_o : n10979_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n10981_o = bf_bset ? n10975_o : n10980_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n10982_o = n10973_o ? n10974_o : n10981_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n10990_o = shifted_bitmask[11];
  /* TG68K_ALU.vhd:592:56  */
  assign n10991_o = result_tmp[11];
  assign n10992_o = n10798_o[11];
  assign n10993_o = n10796_o[11];
  assign n10994_o = n10793_o[11];
  assign n10995_o = n10794_o[11];
  /* TG68K_ALU.vhd:575:17  */
  assign n10996_o = bf_bchg ? n10994_o : n10995_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n10997_o = bf_ins ? n10993_o : n10996_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n10998_o = bf_bset ? n10992_o : n10997_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n10999_o = n10990_o ? n10991_o : n10998_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11007_o = shifted_bitmask[12];
  /* TG68K_ALU.vhd:592:56  */
  assign n11008_o = result_tmp[12];
  assign n11009_o = n10798_o[12];
  assign n11010_o = n10796_o[12];
  assign n11011_o = n10793_o[12];
  assign n11012_o = n10794_o[12];
  /* TG68K_ALU.vhd:575:17  */
  assign n11013_o = bf_bchg ? n11011_o : n11012_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11014_o = bf_ins ? n11010_o : n11013_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11015_o = bf_bset ? n11009_o : n11014_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11016_o = n11007_o ? n11008_o : n11015_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11024_o = shifted_bitmask[13];
  /* TG68K_ALU.vhd:592:56  */
  assign n11025_o = result_tmp[13];
  assign n11026_o = n10798_o[13];
  assign n11027_o = n10796_o[13];
  assign n11028_o = n10793_o[13];
  assign n11029_o = n10794_o[13];
  /* TG68K_ALU.vhd:575:17  */
  assign n11030_o = bf_bchg ? n11028_o : n11029_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11031_o = bf_ins ? n11027_o : n11030_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11032_o = bf_bset ? n11026_o : n11031_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11033_o = n11024_o ? n11025_o : n11032_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11041_o = shifted_bitmask[14];
  /* TG68K_ALU.vhd:592:56  */
  assign n11042_o = result_tmp[14];
  assign n11043_o = n10798_o[14];
  assign n11044_o = n10796_o[14];
  assign n11045_o = n10793_o[14];
  assign n11046_o = n10794_o[14];
  /* TG68K_ALU.vhd:575:17  */
  assign n11047_o = bf_bchg ? n11045_o : n11046_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11048_o = bf_ins ? n11044_o : n11047_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11049_o = bf_bset ? n11043_o : n11048_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11050_o = n11041_o ? n11042_o : n11049_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11058_o = shifted_bitmask[15];
  /* TG68K_ALU.vhd:592:56  */
  assign n11059_o = result_tmp[15];
  assign n11060_o = n10798_o[15];
  assign n11061_o = n10796_o[15];
  assign n11062_o = n10793_o[15];
  assign n11063_o = n10794_o[15];
  /* TG68K_ALU.vhd:575:17  */
  assign n11064_o = bf_bchg ? n11062_o : n11063_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11065_o = bf_ins ? n11061_o : n11064_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11066_o = bf_bset ? n11060_o : n11065_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11067_o = n11058_o ? n11059_o : n11066_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11075_o = shifted_bitmask[16];
  /* TG68K_ALU.vhd:592:56  */
  assign n11076_o = result_tmp[16];
  assign n11077_o = n10798_o[16];
  assign n11078_o = n10796_o[16];
  assign n11079_o = n10793_o[16];
  assign n11080_o = n10794_o[16];
  /* TG68K_ALU.vhd:575:17  */
  assign n11081_o = bf_bchg ? n11079_o : n11080_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11082_o = bf_ins ? n11078_o : n11081_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11083_o = bf_bset ? n11077_o : n11082_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11084_o = n11075_o ? n11076_o : n11083_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11092_o = shifted_bitmask[17];
  /* TG68K_ALU.vhd:592:56  */
  assign n11093_o = result_tmp[17];
  assign n11094_o = n10798_o[17];
  assign n11095_o = n10796_o[17];
  assign n11096_o = n10793_o[17];
  assign n11097_o = n10794_o[17];
  /* TG68K_ALU.vhd:575:17  */
  assign n11098_o = bf_bchg ? n11096_o : n11097_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11099_o = bf_ins ? n11095_o : n11098_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11100_o = bf_bset ? n11094_o : n11099_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11101_o = n11092_o ? n11093_o : n11100_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11109_o = shifted_bitmask[18];
  /* TG68K_ALU.vhd:592:56  */
  assign n11110_o = result_tmp[18];
  assign n11111_o = n10798_o[18];
  assign n11112_o = n10796_o[18];
  assign n11113_o = n10793_o[18];
  assign n11114_o = n10794_o[18];
  /* TG68K_ALU.vhd:575:17  */
  assign n11115_o = bf_bchg ? n11113_o : n11114_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11116_o = bf_ins ? n11112_o : n11115_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11117_o = bf_bset ? n11111_o : n11116_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11118_o = n11109_o ? n11110_o : n11117_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11126_o = shifted_bitmask[19];
  /* TG68K_ALU.vhd:592:56  */
  assign n11127_o = result_tmp[19];
  assign n11128_o = n10798_o[19];
  assign n11129_o = n10796_o[19];
  assign n11130_o = n10793_o[19];
  assign n11131_o = n10794_o[19];
  /* TG68K_ALU.vhd:575:17  */
  assign n11132_o = bf_bchg ? n11130_o : n11131_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11133_o = bf_ins ? n11129_o : n11132_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11134_o = bf_bset ? n11128_o : n11133_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11135_o = n11126_o ? n11127_o : n11134_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11143_o = shifted_bitmask[20];
  /* TG68K_ALU.vhd:592:56  */
  assign n11144_o = result_tmp[20];
  assign n11145_o = n10798_o[20];
  assign n11146_o = n10796_o[20];
  assign n11147_o = n10793_o[20];
  assign n11148_o = n10794_o[20];
  /* TG68K_ALU.vhd:575:17  */
  assign n11149_o = bf_bchg ? n11147_o : n11148_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11150_o = bf_ins ? n11146_o : n11149_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11151_o = bf_bset ? n11145_o : n11150_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11152_o = n11143_o ? n11144_o : n11151_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11160_o = shifted_bitmask[21];
  /* TG68K_ALU.vhd:592:56  */
  assign n11161_o = result_tmp[21];
  assign n11162_o = n10798_o[21];
  assign n11163_o = n10796_o[21];
  assign n11164_o = n10793_o[21];
  assign n11165_o = n10794_o[21];
  /* TG68K_ALU.vhd:575:17  */
  assign n11166_o = bf_bchg ? n11164_o : n11165_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11167_o = bf_ins ? n11163_o : n11166_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11168_o = bf_bset ? n11162_o : n11167_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11169_o = n11160_o ? n11161_o : n11168_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11177_o = shifted_bitmask[22];
  /* TG68K_ALU.vhd:592:56  */
  assign n11178_o = result_tmp[22];
  assign n11179_o = n10798_o[22];
  assign n11180_o = n10796_o[22];
  assign n11181_o = n10793_o[22];
  assign n11182_o = n10794_o[22];
  /* TG68K_ALU.vhd:575:17  */
  assign n11183_o = bf_bchg ? n11181_o : n11182_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11184_o = bf_ins ? n11180_o : n11183_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11185_o = bf_bset ? n11179_o : n11184_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11186_o = n11177_o ? n11178_o : n11185_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11194_o = shifted_bitmask[23];
  /* TG68K_ALU.vhd:592:56  */
  assign n11195_o = result_tmp[23];
  assign n11196_o = n10798_o[23];
  assign n11197_o = n10796_o[23];
  assign n11198_o = n10793_o[23];
  assign n11199_o = n10794_o[23];
  /* TG68K_ALU.vhd:575:17  */
  assign n11200_o = bf_bchg ? n11198_o : n11199_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11201_o = bf_ins ? n11197_o : n11200_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11202_o = bf_bset ? n11196_o : n11201_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11203_o = n11194_o ? n11195_o : n11202_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11211_o = shifted_bitmask[24];
  /* TG68K_ALU.vhd:592:56  */
  assign n11212_o = result_tmp[24];
  assign n11213_o = n10798_o[24];
  assign n11214_o = n10796_o[24];
  assign n11215_o = n10793_o[24];
  assign n11216_o = n10794_o[24];
  /* TG68K_ALU.vhd:575:17  */
  assign n11217_o = bf_bchg ? n11215_o : n11216_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11218_o = bf_ins ? n11214_o : n11217_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11219_o = bf_bset ? n11213_o : n11218_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11220_o = n11211_o ? n11212_o : n11219_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11228_o = shifted_bitmask[25];
  /* TG68K_ALU.vhd:592:56  */
  assign n11229_o = result_tmp[25];
  assign n11230_o = n10798_o[25];
  assign n11231_o = n10796_o[25];
  assign n11232_o = n10793_o[25];
  assign n11233_o = n10794_o[25];
  /* TG68K_ALU.vhd:575:17  */
  assign n11234_o = bf_bchg ? n11232_o : n11233_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11235_o = bf_ins ? n11231_o : n11234_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11236_o = bf_bset ? n11230_o : n11235_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11237_o = n11228_o ? n11229_o : n11236_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11245_o = shifted_bitmask[26];
  /* TG68K_ALU.vhd:592:56  */
  assign n11246_o = result_tmp[26];
  assign n11247_o = n10798_o[26];
  assign n11248_o = n10796_o[26];
  assign n11249_o = n10793_o[26];
  assign n11250_o = n10794_o[26];
  /* TG68K_ALU.vhd:575:17  */
  assign n11251_o = bf_bchg ? n11249_o : n11250_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11252_o = bf_ins ? n11248_o : n11251_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11253_o = bf_bset ? n11247_o : n11252_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11254_o = n11245_o ? n11246_o : n11253_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11262_o = shifted_bitmask[27];
  /* TG68K_ALU.vhd:592:56  */
  assign n11263_o = result_tmp[27];
  assign n11264_o = n10798_o[27];
  assign n11265_o = n10796_o[27];
  assign n11266_o = n10793_o[27];
  assign n11267_o = n10794_o[27];
  /* TG68K_ALU.vhd:575:17  */
  assign n11268_o = bf_bchg ? n11266_o : n11267_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11269_o = bf_ins ? n11265_o : n11268_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11270_o = bf_bset ? n11264_o : n11269_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11271_o = n11262_o ? n11263_o : n11270_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11279_o = shifted_bitmask[28];
  /* TG68K_ALU.vhd:592:56  */
  assign n11280_o = result_tmp[28];
  assign n11281_o = n10798_o[28];
  assign n11282_o = n10796_o[28];
  assign n11283_o = n10793_o[28];
  assign n11284_o = n10794_o[28];
  /* TG68K_ALU.vhd:575:17  */
  assign n11285_o = bf_bchg ? n11283_o : n11284_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11286_o = bf_ins ? n11282_o : n11285_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11287_o = bf_bset ? n11281_o : n11286_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11288_o = n11279_o ? n11280_o : n11287_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11296_o = shifted_bitmask[29];
  /* TG68K_ALU.vhd:592:56  */
  assign n11297_o = result_tmp[29];
  assign n11298_o = n10798_o[29];
  assign n11299_o = n10796_o[29];
  assign n11300_o = n10793_o[29];
  assign n11301_o = n10794_o[29];
  /* TG68K_ALU.vhd:575:17  */
  assign n11302_o = bf_bchg ? n11300_o : n11301_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11303_o = bf_ins ? n11299_o : n11302_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11304_o = bf_bset ? n11298_o : n11303_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11305_o = n11296_o ? n11297_o : n11304_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11313_o = shifted_bitmask[30];
  /* TG68K_ALU.vhd:592:56  */
  assign n11314_o = result_tmp[30];
  assign n11315_o = n10798_o[30];
  assign n11316_o = n10796_o[30];
  assign n11317_o = n10793_o[30];
  assign n11318_o = n10794_o[30];
  /* TG68K_ALU.vhd:575:17  */
  assign n11319_o = bf_bchg ? n11317_o : n11318_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11320_o = bf_ins ? n11316_o : n11319_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11321_o = bf_bset ? n11315_o : n11320_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11322_o = n11313_o ? n11314_o : n11321_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11330_o = shifted_bitmask[31];
  /* TG68K_ALU.vhd:592:56  */
  assign n11331_o = result_tmp[31];
  assign n11332_o = n10798_o[31];
  assign n11333_o = n10796_o[31];
  assign n11334_o = n10793_o[31];
  assign n11335_o = n10794_o[31];
  /* TG68K_ALU.vhd:575:17  */
  assign n11336_o = bf_bchg ? n11334_o : n11335_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11337_o = bf_ins ? n11333_o : n11336_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11338_o = bf_bset ? n11332_o : n11337_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11339_o = n11330_o ? n11331_o : n11338_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11347_o = shifted_bitmask[32];
  /* TG68K_ALU.vhd:592:56  */
  assign n11348_o = result_tmp[32];
  assign n11349_o = n10798_o[32];
  assign n11350_o = n10796_o[32];
  assign n11351_o = n10793_o[32];
  assign n11352_o = n10794_o[32];
  /* TG68K_ALU.vhd:575:17  */
  assign n11353_o = bf_bchg ? n11351_o : n11352_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11354_o = bf_ins ? n11350_o : n11353_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11355_o = bf_bset ? n11349_o : n11354_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11356_o = n11347_o ? n11348_o : n11355_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11364_o = shifted_bitmask[33];
  /* TG68K_ALU.vhd:592:56  */
  assign n11365_o = result_tmp[33];
  assign n11366_o = n10798_o[33];
  assign n11367_o = n10796_o[33];
  assign n11368_o = n10793_o[33];
  assign n11369_o = n10794_o[33];
  /* TG68K_ALU.vhd:575:17  */
  assign n11370_o = bf_bchg ? n11368_o : n11369_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11371_o = bf_ins ? n11367_o : n11370_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11372_o = bf_bset ? n11366_o : n11371_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11373_o = n11364_o ? n11365_o : n11372_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11381_o = shifted_bitmask[34];
  /* TG68K_ALU.vhd:592:56  */
  assign n11382_o = result_tmp[34];
  assign n11383_o = n10798_o[34];
  assign n11384_o = n10796_o[34];
  assign n11385_o = n10793_o[34];
  assign n11386_o = n10794_o[34];
  /* TG68K_ALU.vhd:575:17  */
  assign n11387_o = bf_bchg ? n11385_o : n11386_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11388_o = bf_ins ? n11384_o : n11387_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11389_o = bf_bset ? n11383_o : n11388_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11390_o = n11381_o ? n11382_o : n11389_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11398_o = shifted_bitmask[35];
  /* TG68K_ALU.vhd:592:56  */
  assign n11399_o = result_tmp[35];
  assign n11400_o = n10798_o[35];
  assign n11401_o = n10796_o[35];
  assign n11402_o = n10793_o[35];
  assign n11403_o = n10794_o[35];
  /* TG68K_ALU.vhd:575:17  */
  assign n11404_o = bf_bchg ? n11402_o : n11403_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11405_o = bf_ins ? n11401_o : n11404_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11406_o = bf_bset ? n11400_o : n11405_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11407_o = n11398_o ? n11399_o : n11406_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11415_o = shifted_bitmask[36];
  /* TG68K_ALU.vhd:592:56  */
  assign n11416_o = result_tmp[36];
  assign n11417_o = n10798_o[36];
  assign n11418_o = n10796_o[36];
  assign n11419_o = n10793_o[36];
  assign n11420_o = n10794_o[36];
  /* TG68K_ALU.vhd:575:17  */
  assign n11421_o = bf_bchg ? n11419_o : n11420_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11422_o = bf_ins ? n11418_o : n11421_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11423_o = bf_bset ? n11417_o : n11422_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11424_o = n11415_o ? n11416_o : n11423_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11432_o = shifted_bitmask[37];
  /* TG68K_ALU.vhd:592:56  */
  assign n11433_o = result_tmp[37];
  assign n11434_o = n10798_o[37];
  assign n11435_o = n10796_o[37];
  assign n11436_o = n10793_o[37];
  assign n11437_o = n10794_o[37];
  /* TG68K_ALU.vhd:575:17  */
  assign n11438_o = bf_bchg ? n11436_o : n11437_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11439_o = bf_ins ? n11435_o : n11438_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11440_o = bf_bset ? n11434_o : n11439_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11441_o = n11432_o ? n11433_o : n11440_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11449_o = shifted_bitmask[38];
  /* TG68K_ALU.vhd:592:56  */
  assign n11450_o = result_tmp[38];
  assign n11451_o = n10798_o[38];
  assign n11452_o = n10796_o[38];
  assign n11453_o = n10793_o[38];
  assign n11454_o = n10794_o[38];
  /* TG68K_ALU.vhd:575:17  */
  assign n11455_o = bf_bchg ? n11453_o : n11454_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11456_o = bf_ins ? n11452_o : n11455_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11457_o = bf_bset ? n11451_o : n11456_o;
  /* TG68K_ALU.vhd:591:25  */
  assign n11458_o = n11449_o ? n11450_o : n11457_o;
  assign n11459_o = n10798_o[39];
  assign n11460_o = n10796_o[39];
  assign n11461_o = n10793_o[39];
  assign n11462_o = n10794_o[39];
  /* TG68K_ALU.vhd:575:17  */
  assign n11463_o = bf_bchg ? n11461_o : n11462_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n11464_o = bf_ins ? n11460_o : n11463_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n11465_o = bf_bset ? n11459_o : n11464_o;
  /* TG68K_ALU.vhd:591:43  */
  assign n11466_o = shifted_bitmask[39];
  /* TG68K_ALU.vhd:592:56  */
  assign n11467_o = result_tmp[39];
  /* TG68K_ALU.vhd:591:25  */
  assign n11468_o = n11466_o ? n11467_o : n11465_o;
  /* TG68K_ALU.vhd:598:36  */
  assign n11470_o = {1'b0, bitnr};
  /* TG68K_ALU.vhd:598:43  */
  assign n11471_o = {5'b0, mask_not_zero};  //  uext
  /* TG68K_ALU.vhd:598:43  */
  assign n11472_o = n11470_o + n11471_o;
  /* TG68K_ALU.vhd:601:24  */
  assign n11473_o = mask[31:28];
  /* TG68K_ALU.vhd:601:38  */
  assign n11475_o = n11473_o == 4'b0000;
  /* TG68K_ALU.vhd:602:32  */
  assign n11476_o = mask[27:24];
  /* TG68K_ALU.vhd:602:46  */
  assign n11478_o = n11476_o == 4'b0000;
  /* TG68K_ALU.vhd:603:40  */
  assign n11479_o = mask[23:20];
  /* TG68K_ALU.vhd:603:54  */
  assign n11481_o = n11479_o == 4'b0000;
  /* TG68K_ALU.vhd:604:48  */
  assign n11482_o = mask[19:16];
  /* TG68K_ALU.vhd:604:62  */
  assign n11484_o = n11482_o == 4'b0000;
  /* TG68K_ALU.vhd:606:56  */
  assign n11486_o = mask[15:12];
  /* TG68K_ALU.vhd:606:70  */
  assign n11488_o = n11486_o == 4'b0000;
  /* TG68K_ALU.vhd:607:64  */
  assign n11489_o = mask[11:8];
  /* TG68K_ALU.vhd:607:77  */
  assign n11491_o = n11489_o == 4'b0000;
  /* TG68K_ALU.vhd:609:72  */
  assign n11493_o = mask[7:4];
  /* TG68K_ALU.vhd:609:84  */
  assign n11495_o = n11493_o == 4'b0000;
  /* TG68K_ALU.vhd:611:84  */
  assign n11497_o = mask[3:0];
  /* TG68K_ALU.vhd:613:84  */
  assign n11498_o = mask[7:4];
  /* TG68K_ALU.vhd:609:65  */
  assign n11499_o = n11495_o ? n11497_o : n11498_o;
  /* TG68K_ALU.vhd:609:65  */
  assign n11501_o = n11495_o ? 1'b0 : 1'b1;
  /* TG68K_ALU.vhd:616:76  */
  assign n11502_o = mask[11:8];
  /* TG68K_ALU.vhd:607:57  */
  assign n11504_o = n11491_o ? n11499_o : n11502_o;
  assign n11505_o = {1'b0, n11501_o};
  assign n11506_o = n11505_o[0];
  /* TG68K_ALU.vhd:607:57  */
  assign n11507_o = n11491_o ? n11506_o : 1'b0;
  assign n11508_o = n11505_o[1];
  /* TG68K_ALU.vhd:607:57  */
  assign n11510_o = n11491_o ? n11508_o : 1'b1;
  /* TG68K_ALU.vhd:620:68  */
  assign n11511_o = mask[15:12];
  /* TG68K_ALU.vhd:606:49  */
  assign n11512_o = n11488_o ? n11504_o : n11511_o;
  assign n11513_o = {n11510_o, n11507_o};
  /* TG68K_ALU.vhd:606:49  */
  assign n11515_o = n11488_o ? n11513_o : 2'b11;
  /* TG68K_ALU.vhd:623:60  */
  assign n11516_o = mask[19:16];
  /* TG68K_ALU.vhd:604:41  */
  assign n11519_o = n11484_o ? n11512_o : n11516_o;
  assign n11520_o = {1'b0, 1'b0};
  assign n11521_o = {1'b0, n11515_o};
  assign n11522_o = n11521_o[1:0];
  /* TG68K_ALU.vhd:604:41  */
  assign n11523_o = n11484_o ? n11522_o : n11520_o;
  assign n11524_o = n11521_o[2];
  /* TG68K_ALU.vhd:604:41  */
  assign n11526_o = n11484_o ? n11524_o : 1'b1;
  /* TG68K_ALU.vhd:628:52  */
  assign n11527_o = mask[23:20];
  /* TG68K_ALU.vhd:603:33  */
  assign n11529_o = n11481_o ? n11519_o : n11527_o;
  assign n11530_o = {n11526_o, n11523_o};
  assign n11531_o = n11530_o[0];
  /* TG68K_ALU.vhd:603:33  */
  assign n11533_o = n11481_o ? n11531_o : 1'b1;
  assign n11534_o = n11530_o[1];
  /* TG68K_ALU.vhd:603:33  */
  assign n11535_o = n11481_o ? n11534_o : 1'b0;
  assign n11536_o = n11530_o[2];
  /* TG68K_ALU.vhd:603:33  */
  assign n11538_o = n11481_o ? n11536_o : 1'b1;
  /* TG68K_ALU.vhd:632:44  */
  assign n11539_o = mask[27:24];
  /* TG68K_ALU.vhd:602:25  */
  assign n11541_o = n11478_o ? n11529_o : n11539_o;
  assign n11542_o = {n11538_o, n11535_o, n11533_o};
  assign n11543_o = n11542_o[0];
  /* TG68K_ALU.vhd:602:25  */
  assign n11544_o = n11478_o ? n11543_o : 1'b0;
  assign n11545_o = n11542_o[2:1];
  /* TG68K_ALU.vhd:602:25  */
  assign n11547_o = n11478_o ? n11545_o : 2'b11;
  /* TG68K_ALU.vhd:636:36  */
  assign n11548_o = mask[31:28];
  /* TG68K_ALU.vhd:601:17  */
  assign n11549_o = n11475_o ? n11541_o : n11548_o;
  assign n11550_o = {n11547_o, n11544_o};
  /* TG68K_ALU.vhd:601:17  */
  assign n11552_o = n11475_o ? n11550_o : 3'b111;
  /* TG68K_ALU.vhd:639:23  */
  assign n11555_o = mux[3:2];
  /* TG68K_ALU.vhd:639:35  */
  assign n11557_o = n11555_o == 2'b00;
  /* TG68K_ALU.vhd:641:31  */
  assign n11559_o = mux[1];
  /* TG68K_ALU.vhd:641:34  */
  assign n11560_o = ~n11559_o;
  /* TG68K_ALU.vhd:643:39  */
  assign n11562_o = mux[0];
  /* TG68K_ALU.vhd:643:42  */
  assign n11563_o = ~n11562_o;
  /* TG68K_ALU.vhd:643:33  */
  assign n11566_o = n11563_o ? 1'b0 : 1'b1;
  assign n11567_o = n11553_o[0];
  /* TG68K_ALU.vhd:641:25  */
  assign n11568_o = n11560_o ? 1'b0 : n11567_o;
  /* TG68K_ALU.vhd:641:25  */
  assign n11570_o = n11560_o ? n11566_o : 1'b1;
  /* TG68K_ALU.vhd:648:31  */
  assign n11571_o = mux[3];
  /* TG68K_ALU.vhd:648:34  */
  assign n11572_o = ~n11571_o;
  assign n11574_o = n11553_o[0];
  /* TG68K_ALU.vhd:648:25  */
  assign n11575_o = n11572_o ? 1'b0 : n11574_o;
  assign n11576_o = {1'b0, n11568_o};
  assign n11577_o = n11576_o[0];
  /* TG68K_ALU.vhd:639:17  */
  assign n11578_o = n11557_o ? n11577_o : n11575_o;
  assign n11579_o = n11576_o[1];
  assign n11580_o = n11553_o[1];
  /* TG68K_ALU.vhd:639:17  */
  assign n11581_o = n11557_o ? n11579_o : n11580_o;
  /* TG68K_ALU.vhd:639:17  */
  assign n11584_o = n11557_o ? n11570_o : 1'b1;
  /* TG68K_ALU.vhd:659:32  */
  assign n11589_o = exe_opcode[7:6];
  /* TG68K_ALU.vhd:661:66  */
  assign n11590_o = op1out[7];
  /* TG68K_ALU.vhd:660:25  */
  assign n11592_o = n11589_o == 2'b00;
  /* TG68K_ALU.vhd:663:66  */
  assign n11593_o = op1out[15];
  /* TG68K_ALU.vhd:662:25  */
  assign n11595_o = n11589_o == 2'b01;
  /* TG68K_ALU.vhd:662:34  */
  assign n11597_o = n11589_o == 2'b11;
  /* TG68K_ALU.vhd:662:34  */
  assign n11598_o = n11595_o | n11597_o;
  /* TG68K_ALU.vhd:665:66  */
  assign n11599_o = op1out[31];
  /* TG68K_ALU.vhd:664:25  */
  assign n11601_o = n11589_o == 2'b10;
  assign n11602_o = {n11601_o, n11598_o, n11592_o};
  /* TG68K_ALU.vhd:659:17  */
  always @*
    case (n11602_o)
      3'b100: n11603_o = n11599_o;
      3'b010: n11603_o = n11593_o;
      3'b001: n11603_o = n11590_o;
      default: n11603_o = rot_rot;
    endcase
  /* TG68K_ALU.vhd:670:25  */
  assign n11605_o = rot_bits == 2'b00;
  /* TG68K_ALU.vhd:673:25  */
  assign n11607_o = rot_bits == 2'b01;
  /* TG68K_ALU.vhd:677:65  */
  assign n11608_o = n12821_q[4];
  /* TG68K_ALU.vhd:678:65  */
  assign n11609_o = n12821_q[4];
  /* TG68K_ALU.vhd:676:25  */
  assign n11611_o = rot_bits == 2'b10;
  /* TG68K_ALU.vhd:681:66  */
  assign n11612_o = op1out[0];
  /* TG68K_ALU.vhd:679:25  */
  assign n11614_o = rot_bits == 2'b11;
  assign n11615_o = {n11614_o, n11611_o, n11607_o, n11605_o};
  /* TG68K_ALU.vhd:669:17  */
  always @*
    case (n11615_o)
      4'b1000: n11618_o = rot_rot;
      4'b0100: n11618_o = n11608_o;
      4'b0010: n11618_o = 1'b0;
      4'b0001: n11618_o = 1'b0;
      default: n11618_o = rot_lsb;
    endcase
  /* TG68K_ALU.vhd:669:17  */
  always @*
    case (n11615_o)
      4'b1000: n11620_o = n11612_o;
      4'b0100: n11620_o = n11609_o;
      4'b0010: n11620_o = 1'b0;
      4'b0001: n11620_o = rot_rot;
      default: n11620_o = rot_msb;
    endcase
  /* TG68K_ALU.vhd:685:24  */
  assign n11621_o = exec[23];
  /* TG68K_ALU.vhd:687:39  */
  assign n11622_o = n12821_q[4];
  /* TG68K_ALU.vhd:688:36  */
  assign n11624_o = rot_bits == 2'b10;
  /* TG68K_ALU.vhd:689:47  */
  assign n11625_o = n12821_q[4];
  /* TG68K_ALU.vhd:688:25  */
  assign n11627_o = n11624_o ? n11625_o : 1'b0;
  /* TG68K_ALU.vhd:694:38  */
  assign n11628_o = exe_opcode[8];
  /* TG68K_ALU.vhd:695:50  */
  assign n11629_o = op1out[30:0];
  /* TG68K_ALU.vhd:695:63  */
  assign n11630_o = {n11629_o, rot_lsb};
  /* TG68K_ALU.vhd:699:48  */
  assign n11631_o = op1out[0];
  /* TG68K_ALU.vhd:700:48  */
  assign n11632_o = op1out[0];
  /* TG68K_ALU.vhd:701:58  */
  assign n11633_o = op1out[31:1];
  /* TG68K_ALU.vhd:701:51  */
  assign n11634_o = {rot_msb, n11633_o};
  /* TG68K_ALU.vhd:702:48  */
  assign n11635_o = exe_opcode[7:6];
  /* TG68K_ALU.vhd:703:41  */
  assign n11637_o = n11635_o == 2'b00;
  /* TG68K_ALU.vhd:705:41  */
  assign n11639_o = n11635_o == 2'b01;
  /* TG68K_ALU.vhd:705:50  */
  assign n11641_o = n11635_o == 2'b11;
  /* TG68K_ALU.vhd:705:50  */
  assign n11642_o = n11639_o | n11641_o;
  assign n11643_o = {n11642_o, n11637_o};
  assign n11644_o = n11634_o[7];
  /* TG68K_ALU.vhd:702:33  */
  always @*
    case (n11643_o)
      2'b10: n11645_o = n11644_o;
      2'b01: n11645_o = rot_msb;
      default: n11645_o = n11644_o;
    endcase
  assign n11646_o = n11634_o[15];
  /* TG68K_ALU.vhd:702:33  */
  always @*
    case (n11643_o)
      2'b10: n11647_o = rot_msb;
      2'b01: n11647_o = n11646_o;
      default: n11647_o = n11646_o;
    endcase
  assign n11649_o = n11634_o[6:0];
  assign n11650_o = n11634_o[31:16];
  assign n11651_o = n11634_o[14:8];
  /* TG68K_ALU.vhd:694:25  */
  assign n11652_o = n11628_o ? rot_rot : n11631_o;
  /* TG68K_ALU.vhd:694:25  */
  assign n11653_o = n11628_o ? rot_rot : n11632_o;
  assign n11654_o = {n11650_o, n11647_o, n11651_o, n11645_o, n11649_o};
  /* TG68K_ALU.vhd:694:25  */
  assign n11655_o = n11628_o ? n11630_o : n11654_o;
  /* TG68K_ALU.vhd:685:17  */
  assign n11656_o = n11621_o ? n11622_o : n11652_o;
  /* TG68K_ALU.vhd:685:17  */
  assign n11657_o = n11621_o ? n11627_o : n11653_o;
  /* TG68K_ALU.vhd:685:17  */
  assign n11658_o = n11621_o ? op1out : n11655_o;
  /* TG68K_ALU.vhd:723:28  */
  assign n11663_o = rot_bits == 2'b10;
  /* TG68K_ALU.vhd:724:40  */
  assign n11664_o = exe_opcode[7:6];
  /* TG68K_ALU.vhd:725:33  */
  assign n11666_o = n11664_o == 2'b00;
  /* TG68K_ALU.vhd:727:33  */
  assign n11668_o = n11664_o == 2'b01;
  /* TG68K_ALU.vhd:727:42  */
  assign n11670_o = n11664_o == 2'b11;
  /* TG68K_ALU.vhd:727:42  */
  assign n11671_o = n11668_o | n11670_o;
  /* TG68K_ALU.vhd:729:33  */
  assign n11673_o = n11664_o == 2'b10;
  assign n11674_o = {n11673_o, n11671_o, n11666_o};
  /* TG68K_ALU.vhd:724:25  */
  always @*
    case (n11674_o)
      3'b100: n11679_o = 6'b100001;
      3'b010: n11679_o = 6'b010001;
      3'b001: n11679_o = 6'b001001;
      default: n11679_o = 6'b100000;
    endcase
  /* TG68K_ALU.vhd:734:40  */
  assign n11680_o = exe_opcode[7:6];
  /* TG68K_ALU.vhd:735:33  */
  assign n11682_o = n11680_o == 2'b00;
  /* TG68K_ALU.vhd:737:33  */
  assign n11684_o = n11680_o == 2'b01;
  /* TG68K_ALU.vhd:737:42  */
  assign n11686_o = n11680_o == 2'b11;
  /* TG68K_ALU.vhd:737:42  */
  assign n11687_o = n11684_o | n11686_o;
  /* TG68K_ALU.vhd:739:33  */
  assign n11689_o = n11680_o == 2'b10;
  assign n11690_o = {n11689_o, n11687_o, n11682_o};
  /* TG68K_ALU.vhd:734:25  */
  always @*
    case (n11690_o)
      3'b100: n11695_o = 6'b100000;
      3'b010: n11695_o = 6'b010000;
      3'b001: n11695_o = 6'b001000;
      default: n11695_o = 6'b100000;
    endcase
  /* TG68K_ALU.vhd:723:17  */
  assign n11696_o = n11663_o ? n11679_o : n11695_o;
  /* TG68K_ALU.vhd:745:30  */
  assign n11698_o = exe_opcode[7:6];
  /* TG68K_ALU.vhd:745:42  */
  assign n11700_o = n11698_o == 2'b11;
  /* TG68K_ALU.vhd:745:55  */
  assign n11701_o = exec[81];
  /* TG68K_ALU.vhd:745:64  */
  assign n11702_o = ~n11701_o;
  /* TG68K_ALU.vhd:745:48  */
  assign n11703_o = n11700_o | n11702_o;
  /* TG68K_ALU.vhd:747:33  */
  assign n11704_o = exe_opcode[5];
  /* TG68K_ALU.vhd:748:43  */
  assign n11705_o = op2out[5:0];
  /* TG68K_ALU.vhd:750:59  */
  assign n11706_o = exe_opcode[11:9];
  /* TG68K_ALU.vhd:751:38  */
  assign n11707_o = exe_opcode[11:9];
  /* TG68K_ALU.vhd:751:51  */
  assign n11709_o = n11707_o == 3'b000;
  /* TG68K_ALU.vhd:751:25  */
  assign n11712_o = n11709_o ? 3'b001 : 3'b000;
  assign n11713_o = {n11712_o, n11706_o};
  /* TG68K_ALU.vhd:747:17  */
  assign n11714_o = n11704_o ? n11705_o : n11713_o;
  /* TG68K_ALU.vhd:745:17  */
  assign n11716_o = n11703_o ? 6'b000001 : n11714_o;
  /* TG68K_ALU.vhd:762:29  */
  assign n11723_o = $unsigned(bs_shift) < $unsigned(ring);
  /* TG68K_ALU.vhd:763:40  */
  assign n11724_o = ring - bs_shift;
  /* TG68K_ALU.vhd:762:17  */
  assign n11726_o = n11723_o ? n11724_o : 6'b000000;
  /* TG68K_ALU.vhd:765:45  */
  assign n11728_o = vector[30:0];
  /* TG68K_ALU.vhd:765:38  */
  assign n11730_o = {1'b0, n11728_o};
  /* TG68K_ALU.vhd:765:75  */
  assign n11731_o = vector[31:1];
  /* TG68K_ALU.vhd:765:68  */
  assign n11733_o = {1'b0, n11731_o};
  /* TG68K_ALU.vhd:765:60  */
  assign n11734_o = n11730_o ^ n11733_o;
  /* TG68K_ALU.vhd:765:90  */
  assign n11735_o = {n11734_o, msb};
  /* TG68K_ALU.vhd:766:32  */
  assign n11736_o = exe_opcode[7:6];
  /* TG68K_ALU.vhd:767:25  */
  assign n11739_o = n11736_o == 2'b00;
  /* TG68K_ALU.vhd:769:25  */
  assign n11742_o = n11736_o == 2'b01;
  /* TG68K_ALU.vhd:769:34  */
  assign n11744_o = n11736_o == 2'b11;
  /* TG68K_ALU.vhd:769:34  */
  assign n11745_o = n11742_o | n11744_o;
  assign n11746_o = {n11745_o, n11739_o};
  assign n11747_o = n11735_o[8];
  /* TG68K_ALU.vhd:766:17  */
  always @*
    case (n11746_o)
      2'b10: n11748_o = n11747_o;
      2'b01: n11748_o = 1'b0;
      default: n11748_o = n11747_o;
    endcase
  assign n11749_o = n11735_o[16];
  /* TG68K_ALU.vhd:766:17  */
  always @*
    case (n11746_o)
      2'b10: n11750_o = 1'b0;
      2'b01: n11750_o = n11749_o;
      default: n11750_o = n11749_o;
    endcase
  assign n11752_o = n11735_o[7:0];
  assign n11753_o = n11735_o[32:17];
  assign n11754_o = n11735_o[15:9];
  /* TG68K_ALU.vhd:773:56  */
  assign n11755_o = hot_msb[31:0];
  /* TG68K_ALU.vhd:773:48  */
  assign n11757_o = {1'b0, n11755_o};
  /* TG68K_ALU.vhd:773:42  */
  assign n11758_o = asl_over_xor - n11757_o;
  /* TG68K_ALU.vhd:775:28  */
  assign n11760_o = rot_bits == 2'b00;
  /* TG68K_ALU.vhd:775:48  */
  assign n11761_o = exe_opcode[8];
  /* TG68K_ALU.vhd:775:34  */
  assign n11762_o = n11761_o & n11760_o;
  /* TG68K_ALU.vhd:776:45  */
  assign n11763_o = asl_over[32];
  /* TG68K_ALU.vhd:776:33  */
  assign n11764_o = ~n11763_o;
  /* TG68K_ALU.vhd:775:17  */
  assign n11766_o = n11762_o ? n11764_o : 1'b0;
  /* TG68K_ALU.vhd:780:30  */
  assign n11768_o = exe_opcode[8];
  /* TG68K_ALU.vhd:780:33  */
  assign n11769_o = ~n11768_o;
  /* TG68K_ALU.vhd:781:42  */
  assign n11770_o = result_bs[31];
  /* TG68K_ALU.vhd:783:40  */
  assign n11771_o = exe_opcode[7:6];
  /* TG68K_ALU.vhd:785:58  */
  assign n11772_o = result_bs[8];
  /* TG68K_ALU.vhd:784:33  */
  assign n11774_o = n11771_o == 2'b00;
  /* TG68K_ALU.vhd:787:58  */
  assign n11775_o = result_bs[16];
  /* TG68K_ALU.vhd:786:33  */
  assign n11777_o = n11771_o == 2'b01;
  /* TG68K_ALU.vhd:786:42  */
  assign n11779_o = n11771_o == 2'b11;
  /* TG68K_ALU.vhd:786:42  */
  assign n11780_o = n11777_o | n11779_o;
  /* TG68K_ALU.vhd:789:58  */
  assign n11781_o = result_bs[32];
  /* TG68K_ALU.vhd:788:33  */
  assign n11783_o = n11771_o == 2'b10;
  assign n11784_o = {n11783_o, n11780_o, n11774_o};
  /* TG68K_ALU.vhd:783:25  */
  always @*
    case (n11784_o)
      3'b100: n11785_o = n11781_o;
      3'b010: n11785_o = n11775_o;
      3'b001: n11785_o = n11772_o;
      default: n11785_o = bs_c;
    endcase
  /* TG68K_ALU.vhd:780:17  */
  assign n11786_o = n11769_o ? n11770_o : n11785_o;
  /* TG68K_ALU.vhd:795:28  */
  assign n11788_o = rot_bits == 2'b11;
  /* TG68K_ALU.vhd:796:38  */
  assign n11789_o = n12821_q[4];
  /* TG68K_ALU.vhd:797:40  */
  assign n11790_o = exe_opcode[7:6];
  /* TG68K_ALU.vhd:799:69  */
  assign n11791_o = result_bs[7:0];
  /* TG68K_ALU.vhd:799:94  */
  assign n11792_o = result_bs[15:8];
  /* TG68K_ALU.vhd:799:82  */
  assign n11793_o = n11791_o | n11792_o;
  /* TG68K_ALU.vhd:800:52  */
  assign n11794_o = alu[7];
  /* TG68K_ALU.vhd:798:33  */
  assign n11796_o = n11790_o == 2'b00;
  /* TG68K_ALU.vhd:802:70  */
  assign n11797_o = result_bs[15:0];
  /* TG68K_ALU.vhd:802:96  */
  assign n11798_o = result_bs[31:16];
  /* TG68K_ALU.vhd:802:84  */
  assign n11799_o = n11797_o | n11798_o;
  /* TG68K_ALU.vhd:803:52  */
  assign n11800_o = alu[15];
  /* TG68K_ALU.vhd:801:33  */
  assign n11802_o = n11790_o == 2'b01;
  /* TG68K_ALU.vhd:801:42  */
  assign n11804_o = n11790_o == 2'b11;
  /* TG68K_ALU.vhd:801:42  */
  assign n11805_o = n11802_o | n11804_o;
  /* TG68K_ALU.vhd:805:57  */
  assign n11806_o = result_bs[31:0];
  /* TG68K_ALU.vhd:805:83  */
  assign n11807_o = result_bs[63:32];
  /* TG68K_ALU.vhd:805:71  */
  assign n11808_o = n11806_o | n11807_o;
  /* TG68K_ALU.vhd:806:52  */
  assign n11809_o = alu[31];
  /* TG68K_ALU.vhd:804:33  */
  assign n11811_o = n11790_o == 2'b10;
  assign n11812_o = {n11811_o, n11805_o, n11796_o};
  assign n11813_o = n11799_o[7:0];
  assign n11814_o = n11808_o[7:0];
  /* TG68K_ALU.vhd:797:25  */
  always @*
    case (n11812_o)
      3'b100: n11816_o = n11814_o;
      3'b010: n11816_o = n11813_o;
      3'b001: n11816_o = n11793_o;
      default: n11816_o = 8'bX;
    endcase
  assign n11817_o = n11799_o[15:8];
  assign n11818_o = n11808_o[15:8];
  /* TG68K_ALU.vhd:797:25  */
  always @*
    case (n11812_o)
      3'b100: n11820_o = n11818_o;
      3'b010: n11820_o = n11817_o;
      3'b001: n11820_o = 8'bX;
      default: n11820_o = 8'bX;
    endcase
  assign n11821_o = n11808_o[31:16];
  /* TG68K_ALU.vhd:797:25  */
  always @*
    case (n11812_o)
      3'b100: n11823_o = n11821_o;
      3'b010: n11823_o = 16'bX;
      3'b001: n11823_o = 16'bX;
      default: n11823_o = 16'bX;
    endcase
  /* TG68K_ALU.vhd:797:25  */
  always @*
    case (n11812_o)
      3'b100: n11824_o = n11809_o;
      3'b010: n11824_o = n11800_o;
      3'b001: n11824_o = n11794_o;
      default: n11824_o = n11786_o;
    endcase
  /* TG68K_ALU.vhd:809:38  */
  assign n11825_o = exe_opcode[8];
  /* TG68K_ALU.vhd:810:44  */
  assign n11826_o = alu[0];
  /* TG68K_ALU.vhd:809:25  */
  assign n11827_o = n11825_o ? n11826_o : n11824_o;
  /* TG68K_ALU.vhd:812:31  */
  assign n11829_o = rot_bits == 2'b10;
  /* TG68K_ALU.vhd:813:40  */
  assign n11830_o = exe_opcode[7:6];
  /* TG68K_ALU.vhd:815:69  */
  assign n11831_o = result_bs[7:0];
  /* TG68K_ALU.vhd:815:94  */
  assign n11832_o = result_bs[16:9];
  /* TG68K_ALU.vhd:815:82  */
  assign n11833_o = n11831_o | n11832_o;
  /* TG68K_ALU.vhd:816:58  */
  assign n11834_o = result_bs[8];
  /* TG68K_ALU.vhd:816:74  */
  assign n11835_o = result_bs[17];
  /* TG68K_ALU.vhd:816:62  */
  assign n11836_o = n11834_o | n11835_o;
  /* TG68K_ALU.vhd:814:33  */
  assign n11838_o = n11830_o == 2'b00;
  /* TG68K_ALU.vhd:818:70  */
  assign n11839_o = result_bs[15:0];
  /* TG68K_ALU.vhd:818:96  */
  assign n11840_o = result_bs[32:17];
  /* TG68K_ALU.vhd:818:84  */
  assign n11841_o = n11839_o | n11840_o;
  /* TG68K_ALU.vhd:819:58  */
  assign n11842_o = result_bs[16];
  /* TG68K_ALU.vhd:819:75  */
  assign n11843_o = result_bs[33];
  /* TG68K_ALU.vhd:819:63  */
  assign n11844_o = n11842_o | n11843_o;
  /* TG68K_ALU.vhd:817:33  */
  assign n11846_o = n11830_o == 2'b01;
  /* TG68K_ALU.vhd:817:42  */
  assign n11848_o = n11830_o == 2'b11;
  /* TG68K_ALU.vhd:817:42  */
  assign n11849_o = n11846_o | n11848_o;
  /* TG68K_ALU.vhd:821:57  */
  assign n11850_o = result_bs[31:0];
  /* TG68K_ALU.vhd:821:83  */
  assign n11851_o = result_bs[64:33];
  /* TG68K_ALU.vhd:821:71  */
  assign n11852_o = n11850_o | n11851_o;
  /* TG68K_ALU.vhd:822:58  */
  assign n11853_o = result_bs[32];
  /* TG68K_ALU.vhd:822:75  */
  assign n11854_o = result_bs[65];
  /* TG68K_ALU.vhd:822:63  */
  assign n11855_o = n11853_o | n11854_o;
  /* TG68K_ALU.vhd:820:33  */
  assign n11857_o = n11830_o == 2'b10;
  assign n11858_o = {n11857_o, n11849_o, n11838_o};
  assign n11859_o = n11841_o[7:0];
  assign n11860_o = n11852_o[7:0];
  /* TG68K_ALU.vhd:813:25  */
  always @*
    case (n11858_o)
      3'b100: n11862_o = n11860_o;
      3'b010: n11862_o = n11859_o;
      3'b001: n11862_o = n11833_o;
      default: n11862_o = 8'bX;
    endcase
  assign n11863_o = n11841_o[15:8];
  assign n11864_o = n11852_o[15:8];
  /* TG68K_ALU.vhd:813:25  */
  always @*
    case (n11858_o)
      3'b100: n11866_o = n11864_o;
      3'b010: n11866_o = n11863_o;
      3'b001: n11866_o = 8'bX;
      default: n11866_o = 8'bX;
    endcase
  assign n11867_o = n11852_o[31:16];
  /* TG68K_ALU.vhd:813:25  */
  always @*
    case (n11858_o)
      3'b100: n11869_o = n11867_o;
      3'b010: n11869_o = 16'bX;
      3'b001: n11869_o = 16'bX;
      default: n11869_o = 16'bX;
    endcase
  /* TG68K_ALU.vhd:813:25  */
  always @*
    case (n11858_o)
      3'b100: n11870_o = n11855_o;
      3'b010: n11870_o = n11844_o;
      3'b001: n11870_o = n11836_o;
      default: n11870_o = n11786_o;
    endcase
  /* TG68K_ALU.vhd:826:38  */
  assign n11871_o = exe_opcode[8];
  /* TG68K_ALU.vhd:826:41  */
  assign n11872_o = ~n11871_o;
  /* TG68K_ALU.vhd:827:49  */
  assign n11873_o = result_bs[63:32];
  /* TG68K_ALU.vhd:829:49  */
  assign n11874_o = result_bs[31:0];
  /* TG68K_ALU.vhd:826:25  */
  assign n11875_o = n11872_o ? n11873_o : n11874_o;
  assign n11876_o = {n11869_o, n11866_o, n11862_o};
  /* TG68K_ALU.vhd:812:17  */
  assign n11877_o = n11829_o ? n11876_o : n11875_o;
  /* TG68K_ALU.vhd:812:17  */
  assign n11878_o = n11829_o ? n11870_o : n11786_o;
  assign n11879_o = {n11823_o, n11820_o, n11816_o};
  /* TG68K_ALU.vhd:795:17  */
  assign n11880_o = n11788_o ? n11879_o : n11877_o;
  /* TG68K_ALU.vhd:795:17  */
  assign n11882_o = n11788_o ? n11827_o : n11878_o;
  /* TG68K_ALU.vhd:795:17  */
  assign n11883_o = n11788_o ? n11789_o : bs_c;
  /* TG68K_ALU.vhd:833:29  */
  assign n11885_o = bs_shift == 6'b000000;
  /* TG68K_ALU.vhd:834:36  */
  assign n11887_o = rot_bits == 2'b10;
  /* TG68K_ALU.vhd:835:46  */
  assign n11888_o = n12821_q[4];
  /* TG68K_ALU.vhd:834:25  */
  assign n11890_o = n11887_o ? n11888_o : 1'b0;
  /* TG68K_ALU.vhd:839:38  */
  assign n11891_o = n12821_q[4];
  /* TG68K_ALU.vhd:833:17  */
  assign n11893_o = n11885_o ? 1'b0 : n11766_o;
  /* TG68K_ALU.vhd:833:17  */
  assign n11894_o = n11885_o ? n11890_o : n11882_o;
  /* TG68K_ALU.vhd:833:17  */
  assign n11895_o = n11885_o ? n11891_o : n11883_o;
  /* TG68K_ALU.vhd:848:45  */
  assign n11897_o = bs_shift == 6'b111111;
  /* TG68K_ALU.vhd:850:48  */
  assign n11899_o = $unsigned(bs_shift) > $unsigned(6'b110101);
  /* TG68K_ALU.vhd:851:66  */
  assign n11901_o = bs_shift - 6'b110110;
  /* TG68K_ALU.vhd:852:48  */
  assign n11903_o = $unsigned(bs_shift) > $unsigned(6'b101100);
  /* TG68K_ALU.vhd:853:66  */
  assign n11905_o = bs_shift - 6'b101101;
  /* TG68K_ALU.vhd:854:48  */
  assign n11907_o = $unsigned(bs_shift) > $unsigned(6'b100011);
  /* TG68K_ALU.vhd:855:66  */
  assign n11909_o = bs_shift - 6'b100100;
  /* TG68K_ALU.vhd:856:48  */
  assign n11911_o = $unsigned(bs_shift) > $unsigned(6'b011010);
  /* TG68K_ALU.vhd:857:66  */
  assign n11913_o = bs_shift - 6'b011011;
  /* TG68K_ALU.vhd:858:48  */
  assign n11915_o = $unsigned(bs_shift) > $unsigned(6'b010001);
  /* TG68K_ALU.vhd:859:66  */
  assign n11917_o = bs_shift - 6'b010010;
  /* TG68K_ALU.vhd:860:48  */
  assign n11919_o = $unsigned(bs_shift) > $unsigned(6'b001000);
  /* TG68K_ALU.vhd:861:66  */
  assign n11921_o = bs_shift - 6'b001001;
  /* TG68K_ALU.vhd:860:33  */
  assign n11922_o = n11919_o ? n11921_o : bs_shift;
  /* TG68K_ALU.vhd:858:33  */
  assign n11923_o = n11915_o ? n11917_o : n11922_o;
  /* TG68K_ALU.vhd:856:33  */
  assign n11924_o = n11911_o ? n11913_o : n11923_o;
  /* TG68K_ALU.vhd:854:33  */
  assign n11925_o = n11907_o ? n11909_o : n11924_o;
  /* TG68K_ALU.vhd:852:33  */
  assign n11926_o = n11903_o ? n11905_o : n11925_o;
  /* TG68K_ALU.vhd:850:33  */
  assign n11927_o = n11899_o ? n11901_o : n11926_o;
  /* TG68K_ALU.vhd:848:33  */
  assign n11929_o = n11897_o ? 6'b000000 : n11927_o;
  /* TG68K_ALU.vhd:847:25  */
  assign n11931_o = ring == 6'b001001;
  /* TG68K_ALU.vhd:866:45  */
  assign n11933_o = $unsigned(bs_shift) > $unsigned(6'b110010);
  /* TG68K_ALU.vhd:867:66  */
  assign n11935_o = bs_shift - 6'b110011;
  /* TG68K_ALU.vhd:868:48  */
  assign n11937_o = $unsigned(bs_shift) > $unsigned(6'b100001);
  /* TG68K_ALU.vhd:869:66  */
  assign n11939_o = bs_shift - 6'b100010;
  /* TG68K_ALU.vhd:870:48  */
  assign n11941_o = $unsigned(bs_shift) > $unsigned(6'b010000);
  /* TG68K_ALU.vhd:871:66  */
  assign n11943_o = bs_shift - 6'b010001;
  /* TG68K_ALU.vhd:870:33  */
  assign n11944_o = n11941_o ? n11943_o : bs_shift;
  /* TG68K_ALU.vhd:868:33  */
  assign n11945_o = n11937_o ? n11939_o : n11944_o;
  /* TG68K_ALU.vhd:866:33  */
  assign n11946_o = n11933_o ? n11935_o : n11945_o;
  /* TG68K_ALU.vhd:865:25  */
  assign n11948_o = ring == 6'b010001;
  /* TG68K_ALU.vhd:876:45  */
  assign n11950_o = $unsigned(bs_shift) > $unsigned(6'b100000);
  /* TG68K_ALU.vhd:877:66  */
  assign n11952_o = bs_shift - 6'b100001;
  /* TG68K_ALU.vhd:876:33  */
  assign n11953_o = n11950_o ? n11952_o : bs_shift;
  /* TG68K_ALU.vhd:875:25  */
  assign n11955_o = ring == 6'b100001;
  /* TG68K_ALU.vhd:881:74  */
  assign n11956_o = bs_shift[2:0];
  /* TG68K_ALU.vhd:881:64  */
  assign n11958_o = {3'b000, n11956_o};
  /* TG68K_ALU.vhd:881:25  */
  assign n11960_o = ring == 6'b001000;
  /* TG68K_ALU.vhd:882:74  */
  assign n11961_o = bs_shift[3:0];
  /* TG68K_ALU.vhd:882:64  */
  assign n11963_o = {2'b00, n11961_o};
  /* TG68K_ALU.vhd:882:25  */
  assign n11965_o = ring == 6'b010000;
  /* TG68K_ALU.vhd:883:74  */
  assign n11966_o = bs_shift[4:0];
  /* TG68K_ALU.vhd:883:64  */
  assign n11968_o = {1'b0, n11966_o};
  /* TG68K_ALU.vhd:883:25  */
  assign n11970_o = ring == 6'b100000;
  assign n11971_o = {n11970_o, n11965_o, n11960_o, n11955_o, n11948_o, n11931_o};
  /* TG68K_ALU.vhd:846:17  */
  always @*
    case (n11971_o)
      6'b100000: n11973_o = n11968_o;
      6'b010000: n11973_o = n11963_o;
      6'b001000: n11973_o = n11958_o;
      6'b000100: n11973_o = n11953_o;
      6'b000010: n11973_o = n11946_o;
      6'b000001: n11973_o = n11929_o;
      default: n11973_o = 6'b000000;
    endcase
  /* TG68K_ALU.vhd:888:30  */
  assign n11974_o = exe_opcode[8];
  /* TG68K_ALU.vhd:888:33  */
  assign n11975_o = ~n11974_o;
  /* TG68K_ALU.vhd:889:39  */
  assign n11976_o = ring - bs_shift_mod;
  /* TG68K_ALU.vhd:888:17  */
  assign n11977_o = n11975_o ? n11976_o : bs_shift_mod;
  /* TG68K_ALU.vhd:891:28  */
  assign n11978_o = rot_bits[1];
  /* TG68K_ALU.vhd:891:31  */
  assign n11979_o = ~n11978_o;
  /* TG68K_ALU.vhd:892:38  */
  assign n11980_o = exe_opcode[8];
  /* TG68K_ALU.vhd:892:41  */
  assign n11981_o = ~n11980_o;
  /* TG68K_ALU.vhd:893:45  */
  assign n11983_o = 6'b100000 - bs_shift_mod;
  /* TG68K_ALU.vhd:892:25  */
  assign n11984_o = n11981_o ? n11983_o : n11977_o;
  /* TG68K_ALU.vhd:895:37  */
  assign n11985_o = bs_shift == ring;
  /* TG68K_ALU.vhd:896:46  */
  assign n11986_o = exe_opcode[8];
  /* TG68K_ALU.vhd:896:49  */
  assign n11987_o = ~n11986_o;
  /* TG68K_ALU.vhd:897:53  */
  assign n11989_o = 6'b100000 - ring;
  /* TG68K_ALU.vhd:896:33  */
  assign n11990_o = n11987_o ? n11989_o : ring;
  /* TG68K_ALU.vhd:895:25  */
  assign n11991_o = n11985_o ? n11990_o : n11984_o;
  /* TG68K_ALU.vhd:902:37  */
  assign n11992_o = $unsigned(bs_shift) > $unsigned(ring);
  /* TG68K_ALU.vhd:903:46  */
  assign n11993_o = exe_opcode[8];
  /* TG68K_ALU.vhd:903:49  */
  assign n11994_o = ~n11993_o;
  /* TG68K_ALU.vhd:907:55  */
  assign n11996_o = ring + 6'b000001;
  /* TG68K_ALU.vhd:903:33  */
  assign n11998_o = n11994_o ? 6'b000000 : n11996_o;
  /* TG68K_ALU.vhd:891:17  */
  assign n12000_o = n12004_o ? 1'b0 : n11894_o;
  /* TG68K_ALU.vhd:902:25  */
  assign n12001_o = n11992_o ? n11998_o : n11991_o;
  /* TG68K_ALU.vhd:902:25  */
  assign n12002_o = n11994_o & n11992_o;
  /* TG68K_ALU.vhd:891:17  */
  assign n12003_o = n11979_o ? n12001_o : n11977_o;
  /* TG68K_ALU.vhd:891:17  */
  assign n12004_o = n12002_o & n11979_o;
  /* TG68K_ALU.vhd:915:50  */
  assign n12005_o = asr_sign[31:0];
  /* TG68K_ALU.vhd:915:74  */
  assign n12006_o = hot_msb[31:0];
  /* TG68K_ALU.vhd:915:64  */
  assign n12007_o = n12005_o | n12006_o;
  assign n12009_o = n12008_o[0];
  /* TG68K_ALU.vhd:916:28  */
  assign n12011_o = rot_bits == 2'b00;
  /* TG68K_ALU.vhd:916:48  */
  assign n12012_o = exe_opcode[8];
  /* TG68K_ALU.vhd:916:51  */
  assign n12013_o = ~n12012_o;
  /* TG68K_ALU.vhd:916:34  */
  assign n12014_o = n12013_o & n12011_o;
  /* TG68K_ALU.vhd:916:56  */
  assign n12015_o = msb & n12014_o;
  /* TG68K_ALU.vhd:917:49  */
  assign n12016_o = asr_sign[32:1];
  /* TG68K_ALU.vhd:917:38  */
  assign n12017_o = alu | n12016_o;
  /* TG68K_ALU.vhd:918:37  */
  assign n12018_o = $unsigned(bs_shift) > $unsigned(ring);
  /* TG68K_ALU.vhd:916:17  */
  assign n12020_o = n12022_o ? 1'b1 : n12000_o;
  /* TG68K_ALU.vhd:916:17  */
  assign n12022_o = n12018_o & n12015_o;
  /* TG68K_ALU.vhd:923:43  */
  assign n12024_o = {1'b0, op1out};
  /* TG68K_ALU.vhd:924:32  */
  assign n12025_o = exe_opcode[7:6];
  /* TG68K_ALU.vhd:926:46  */
  assign n12026_o = op1out[7];
  /* TG68K_ALU.vhd:929:44  */
  assign n12030_o = rot_bits == 2'b10;
  /* TG68K_ALU.vhd:930:59  */
  assign n12031_o = n12821_q[4];
  assign n12032_o = n12027_o[0];
  /* TG68K_ALU.vhd:929:33  */
  assign n12033_o = n12030_o ? n12031_o : n12032_o;
  assign n12034_o = n12027_o[23:1];
  /* TG68K_ALU.vhd:925:25  */
  assign n12036_o = n12025_o == 2'b00;
  /* TG68K_ALU.vhd:933:46  */
  assign n12037_o = op1out[15];
  /* TG68K_ALU.vhd:936:44  */
  assign n12041_o = rot_bits == 2'b10;
  /* TG68K_ALU.vhd:937:60  */
  assign n12042_o = n12821_q[4];
  assign n12043_o = n12038_o[0];
  /* TG68K_ALU.vhd:936:33  */
  assign n12044_o = n12041_o ? n12042_o : n12043_o;
  assign n12045_o = n12038_o[15:1];
  /* TG68K_ALU.vhd:932:25  */
  assign n12047_o = n12025_o == 2'b01;
  /* TG68K_ALU.vhd:932:34  */
  assign n12049_o = n12025_o == 2'b11;
  /* TG68K_ALU.vhd:932:34  */
  assign n12050_o = n12047_o | n12049_o;
  /* TG68K_ALU.vhd:940:46  */
  assign n12051_o = op1out[31];
  /* TG68K_ALU.vhd:941:44  */
  assign n12053_o = rot_bits == 2'b10;
  /* TG68K_ALU.vhd:942:60  */
  assign n12054_o = n12821_q[4];
  assign n12055_o = n12024_o[32];
  /* TG68K_ALU.vhd:941:33  */
  assign n12056_o = n12053_o ? n12054_o : n12055_o;
  /* TG68K_ALU.vhd:939:25  */
  assign n12058_o = n12025_o == 2'b10;
  assign n12059_o = {n12058_o, n12050_o, n12036_o};
  assign n12060_o = n12024_o[8];
  /* TG68K_ALU.vhd:924:17  */
  always @*
    case (n12059_o)
      3'b100: n12061_o = n12060_o;
      3'b010: n12061_o = n12060_o;
      3'b001: n12061_o = n12033_o;
      default: n12061_o = n12060_o;
    endcase
  assign n12062_o = n12034_o[6:0];
  assign n12063_o = n12024_o[15:9];
  /* TG68K_ALU.vhd:924:17  */
  always @*
    case (n12059_o)
      3'b100: n12064_o = n12063_o;
      3'b010: n12064_o = n12063_o;
      3'b001: n12064_o = n12062_o;
      default: n12064_o = n12063_o;
    endcase
  assign n12065_o = n12034_o[7];
  assign n12066_o = n12024_o[16];
  /* TG68K_ALU.vhd:924:17  */
  always @*
    case (n12059_o)
      3'b100: n12067_o = n12066_o;
      3'b010: n12067_o = n12044_o;
      3'b001: n12067_o = n12065_o;
      default: n12067_o = n12066_o;
    endcase
  assign n12068_o = n12034_o[22:8];
  assign n12069_o = n12024_o[31:17];
  /* TG68K_ALU.vhd:924:17  */
  always @*
    case (n12059_o)
      3'b100: n12070_o = n12069_o;
      3'b010: n12070_o = n12045_o;
      3'b001: n12070_o = n12068_o;
      default: n12070_o = n12069_o;
    endcase
  assign n12071_o = n12024_o[32];
  /* TG68K_ALU.vhd:924:17  */
  always @*
    case (n12059_o)
      3'b100: n12072_o = n12056_o;
      3'b010: n12072_o = n12071_o;
      3'b001: n12072_o = n12071_o;
      default: n12072_o = n12071_o;
    endcase
  assign n12074_o = n12024_o[7:0];
  /* TG68K_ALU.vhd:924:17  */
  always @*
    case (n12059_o)
      3'b100: n12078_o = n12051_o;
      3'b010: n12078_o = n12037_o;
      3'b001: n12078_o = n12026_o;
      default: n12078_o = msb;
    endcase
  assign n12079_o = n12028_o[7:0];
  assign n12080_o = n12017_o[15:8];
  assign n12081_o = alu[15:8];
  /* TG68K_ALU.vhd:916:17  */
  assign n12082_o = n12015_o ? n12080_o : n12081_o;
  /* TG68K_ALU.vhd:924:17  */
  always @*
    case (n12059_o)
      3'b100: n12083_o = n12082_o;
      3'b010: n12083_o = n12082_o;
      3'b001: n12083_o = n12079_o;
      default: n12083_o = n12082_o;
    endcase
  assign n12084_o = n12028_o[23:8];
  assign n12085_o = n12017_o[31:16];
  assign n12086_o = alu[31:16];
  /* TG68K_ALU.vhd:916:17  */
  assign n12087_o = n12015_o ? n12085_o : n12086_o;
  /* TG68K_ALU.vhd:924:17  */
  always @*
    case (n12059_o)
      3'b100: n12088_o = n12087_o;
      3'b010: n12088_o = 16'b0000000000000000;
      3'b001: n12088_o = n12084_o;
      default: n12088_o = n12087_o;
    endcase
  assign n12092_o = n12017_o[7:0];
  assign n12093_o = alu[7:0];
  /* TG68K_ALU.vhd:916:17  */
  assign n12094_o = n12015_o ? n12092_o : n12093_o;
  /* TG68K_ALU.vhd:946:71  */
  assign n12096_o = {33'b000000000000000000000000000000000, vector};
  /* TG68K_ALU.vhd:946:84  */
  assign n12097_o = {25'b0, bit_nr};  //  uext
  /* TG68K_ALU.vhd:946:80  */
  assign n12098_o = {1'b0, n12097_o};  //  uext
  /* TG68K_ALU.vhd:946:80  */
  assign n12099_o = n12096_o << n12098_o;
  /* TG68K_ALU.vhd:957:24  */
  assign n12103_o = exec[17];
  /* TG68K_ALU.vhd:958:58  */
  assign n12104_o = last_data_read[7:0];
  /* TG68K_ALU.vhd:958:40  */
  assign n12105_o = n12821_q & n12104_o;
  /* TG68K_ALU.vhd:959:27  */
  assign n12106_o = exec[18];
  /* TG68K_ALU.vhd:960:58  */
  assign n12107_o = last_data_read[7:0];
  /* TG68K_ALU.vhd:960:40  */
  assign n12108_o = n12821_q ^ n12107_o;
  /* TG68K_ALU.vhd:961:27  */
  assign n12109_o = exec[19];
  /* TG68K_ALU.vhd:962:57  */
  assign n12110_o = last_data_read[7:0];
  /* TG68K_ALU.vhd:962:40  */
  assign n12111_o = n12821_q | n12110_o;
  /* TG68K_ALU.vhd:964:40  */
  assign n12112_o = op2out[7:0];
  /* TG68K_ALU.vhd:961:17  */
  assign n12113_o = n12109_o ? n12111_o : n12112_o;
  /* TG68K_ALU.vhd:959:17  */
  assign n12114_o = n12106_o ? n12108_o : n12113_o;
  /* TG68K_ALU.vhd:957:17  */
  assign n12115_o = n12103_o ? n12105_o : n12114_o;
  /* TG68K_ALU.vhd:971:24  */
  assign n12116_o = exec[28];
  /* TG68K_ALU.vhd:971:50  */
  assign n12117_o = n12821_q[2];
  /* TG68K_ALU.vhd:971:53  */
  assign n12118_o = ~n12117_o;
  /* TG68K_ALU.vhd:971:41  */
  assign n12119_o = n12118_o & n12116_o;
  /* TG68K_ALU.vhd:973:28  */
  assign n12120_o = op1in[7:0];
  /* TG68K_ALU.vhd:973:40  */
  assign n12122_o = n12120_o == 8'b00000000;
  /* TG68K_ALU.vhd:975:33  */
  assign n12124_o = op1in[15:8];
  /* TG68K_ALU.vhd:975:46  */
  assign n12126_o = n12124_o == 8'b00000000;
  /* TG68K_ALU.vhd:977:41  */
  assign n12128_o = op1in[31:16];
  /* TG68K_ALU.vhd:977:55  */
  assign n12130_o = n12128_o == 16'b0000000000000000;
  /* TG68K_ALU.vhd:977:33  */
  assign n12133_o = n12130_o ? 1'b1 : 1'b0;
  assign n12134_o = {n12133_o, 1'b1};
  /* TG68K_ALU.vhd:975:25  */
  assign n12136_o = n12126_o ? n12134_o : 2'b00;
  assign n12137_o = {n12136_o, 1'b1};
  /* TG68K_ALU.vhd:973:17  */
  assign n12139_o = n12122_o ? n12137_o : 3'b000;
  /* TG68K_ALU.vhd:971:17  */
  assign n12141_o = n12119_o ? 3'b000 : n12139_o;
  /* TG68K_ALU.vhd:984:32  */
  assign n12144_o = exe_datatype == 2'b00;
  /* TG68K_ALU.vhd:985:43  */
  assign n12145_o = op1in[7];
  /* TG68K_ALU.vhd:985:53  */
  assign n12146_o = flag_z[0];
  /* TG68K_ALU.vhd:985:46  */
  assign n12147_o = {n12145_o, n12146_o};
  /* TG68K_ALU.vhd:985:67  */
  assign n12148_o = addsub_ofl[0];
  /* TG68K_ALU.vhd:985:56  */
  assign n12149_o = {n12147_o, n12148_o};
  /* TG68K_ALU.vhd:985:76  */
  assign n12150_o = n10046_o[0];
  /* TG68K_ALU.vhd:985:70  */
  assign n12151_o = {n12149_o, n12150_o};
  /* TG68K_ALU.vhd:986:32  */
  assign n12152_o = exec[12];
  /* TG68K_ALU.vhd:986:53  */
  assign n12153_o = exec[13];
  /* TG68K_ALU.vhd:986:46  */
  assign n12154_o = n12152_o | n12153_o;
  assign n12155_o = {vflag_a, bcd_a_carry};
  assign n12156_o = n12151_o[1:0];
  /* TG68K_ALU.vhd:986:25  */
  assign n12157_o = n12154_o ? n12155_o : n12156_o;
  assign n12158_o = n12151_o[3:2];
  /* TG68K_ALU.vhd:990:35  */
  assign n12160_o = exe_datatype == 2'b10;
  /* TG68K_ALU.vhd:990:48  */
  assign n12161_o = exec[10];
  /* TG68K_ALU.vhd:990:41  */
  assign n12162_o = n12160_o | n12161_o;
  /* TG68K_ALU.vhd:991:43  */
  assign n12163_o = op1in[31];
  /* TG68K_ALU.vhd:991:54  */
  assign n12164_o = flag_z[2];
  /* TG68K_ALU.vhd:991:47  */
  assign n12165_o = {n12163_o, n12164_o};
  /* TG68K_ALU.vhd:991:68  */
  assign n12166_o = addsub_ofl[2];
  /* TG68K_ALU.vhd:991:57  */
  assign n12167_o = {n12165_o, n12166_o};
  /* TG68K_ALU.vhd:991:77  */
  assign n12168_o = n10046_o[2];
  /* TG68K_ALU.vhd:991:71  */
  assign n12169_o = {n12167_o, n12168_o};
  /* TG68K_ALU.vhd:993:43  */
  assign n12170_o = op1in[15];
  /* TG68K_ALU.vhd:993:54  */
  assign n12171_o = flag_z[1];
  /* TG68K_ALU.vhd:993:47  */
  assign n12172_o = {n12170_o, n12171_o};
  /* TG68K_ALU.vhd:993:68  */
  assign n12173_o = addsub_ofl[1];
  /* TG68K_ALU.vhd:993:57  */
  assign n12174_o = {n12172_o, n12173_o};
  /* TG68K_ALU.vhd:993:77  */
  assign n12175_o = n10046_o[1];
  /* TG68K_ALU.vhd:993:71  */
  assign n12176_o = {n12174_o, n12175_o};
  /* TG68K_ALU.vhd:990:17  */
  assign n12177_o = n12162_o ? n12169_o : n12176_o;
  assign n12178_o = {n12158_o, n12157_o};
  /* TG68K_ALU.vhd:984:17  */
  assign n12179_o = n12144_o ? n12178_o : n12177_o;
  /* TG68K_ALU.vhd:1000:40  */
  assign n12181_o = exec[59];
  /* TG68K_ALU.vhd:1000:55  */
  assign n12182_o = n12181_o | set_stop;
  /* TG68K_ALU.vhd:1003:40  */
  assign n12185_o = exec[60];
  /* TG68K_ALU.vhd:1007:40  */
  assign n12188_o = exec[9];
  /* TG68K_ALU.vhd:1007:66  */
  assign n12189_o = ~decodeopc;
  /* TG68K_ALU.vhd:1007:53  */
  assign n12190_o = n12189_o & n12188_o;
  /* TG68K_ALU.vhd:1008:65  */
  assign n12191_o = set_flags[3];
  /* TG68K_ALU.vhd:1008:69  */
  assign n12192_o = n12191_o ^ rot_rot;
  /* TG68K_ALU.vhd:1008:82  */
  assign n12193_o = n12192_o | asl_vflag;
  /* TG68K_ALU.vhd:1007:33  */
  assign n12195_o = n12190_o ? n12193_o : 1'b0;
  /* TG68K_ALU.vhd:1012:40  */
  assign n12196_o = exec[51];
  /* TG68K_ALU.vhd:1015:56  */
  assign n12198_o = micro_state == 7'b0110011;
  /* TG68K_ALU.vhd:1017:62  */
  assign n12199_o = exe_opcode[8];
  /* TG68K_ALU.vhd:1017:65  */
  assign n12200_o = ~n12199_o;
  /* TG68K_ALU.vhd:1019:92  */
  assign n12201_o = reg_qa[31];
  /* TG68K_ALU.vhd:1019:82  */
  assign n12202_o = ~n12201_o;
  /* TG68K_ALU.vhd:1019:81  */
  assign n12204_o = {1'b0, n12202_o};
  /* TG68K_ALU.vhd:1019:96  */
  assign n12206_o = {n12204_o, 2'b00};
  /* TG68K_ALU.vhd:1017:49  */
  assign n12208_o = n12200_o ? n12206_o : 4'b0100;
  assign n12209_o = data_read[3:0];
  assign n12210_o = data_read[3:0];
  assign n12211_o = n12821_q[3:0];
  /* TG68K_ALU.vhd:1000:33  */
  assign n12212_o = n12182_o ? n12210_o : n12211_o;
  /* TG68K_ALU.vhd:1003:33  */
  assign n12213_o = n12185_o ? n12209_o : n12212_o;
  /* TG68K_ALU.vhd:1015:41  */
  assign n12214_o = n12198_o ? n12208_o : n12213_o;
  /* TG68K_ALU.vhd:1024:43  */
  assign n12215_o = exec[49];
  /* TG68K_ALU.vhd:1024:53  */
  assign n12216_o = ~n12215_o;
  /* TG68K_ALU.vhd:1025:61  */
  assign n12217_o = n12821_q[3:0];
  /* TG68K_ALU.vhd:1026:48  */
  assign n12218_o = exec[3];
  /* TG68K_ALU.vhd:1027:70  */
  assign n12219_o = set_flags[0];
  /* TG68K_ALU.vhd:1028:51  */
  assign n12220_o = exec[9];
  /* TG68K_ALU.vhd:1028:76  */
  assign n12222_o = rot_bits != 2'b11;
  /* TG68K_ALU.vhd:1028:64  */
  assign n12223_o = n12222_o & n12220_o;
  /* TG68K_ALU.vhd:1028:91  */
  assign n12224_o = exec[23];
  /* TG68K_ALU.vhd:1028:100  */
  assign n12225_o = ~n12224_o;
  /* TG68K_ALU.vhd:1028:83  */
  assign n12226_o = n12225_o & n12223_o;
  /* TG68K_ALU.vhd:1030:51  */
  assign n12227_o = exec[81];
  assign n12228_o = data_read[4];
  assign n12229_o = data_read[4];
  assign n12230_o = n12821_q[4];
  /* TG68K_ALU.vhd:1000:33  */
  assign n12231_o = n12182_o ? n12229_o : n12230_o;
  /* TG68K_ALU.vhd:1003:33  */
  assign n12232_o = n12185_o ? n12228_o : n12231_o;
  /* TG68K_ALU.vhd:1030:41  */
  assign n12233_o = n12227_o ? bs_x : n12232_o;
  /* TG68K_ALU.vhd:1028:41  */
  assign n12234_o = n12226_o ? rot_x : n12233_o;
  /* TG68K_ALU.vhd:1026:41  */
  assign n12235_o = n12218_o ? n12219_o : n12234_o;
  /* TG68K_ALU.vhd:1034:49  */
  assign n12236_o = exec[8];
  /* TG68K_ALU.vhd:1034:65  */
  assign n12237_o = exec[86];
  /* TG68K_ALU.vhd:1034:58  */
  assign n12238_o = n12236_o | n12237_o;
  /* TG68K_ALU.vhd:1036:51  */
  assign n12239_o = exec[21];
  /* TG68K_ALU.vhd:1036:65  */
  assign n12241_o = 1'b1 & n12239_o;
  /* TG68K_ALU.vhd:1039:65  */
  assign n12243_o = exe_opcode[15];
  /* TG68K_ALU.vhd:1039:74  */
  assign n12245_o = n12243_o | 1'b0;
  /* TG68K_ALU.vhd:1040:83  */
  assign n12246_o = op1in[15];
  /* TG68K_ALU.vhd:1040:94  */
  assign n12247_o = flag_z[1];
  /* TG68K_ALU.vhd:1040:87  */
  assign n12248_o = {n12246_o, n12247_o};
  /* TG68K_ALU.vhd:1040:97  */
  assign n12250_o = {n12248_o, 2'b00};
  /* TG68K_ALU.vhd:1042:83  */
  assign n12251_o = op1in[31];
  /* TG68K_ALU.vhd:1042:94  */
  assign n12252_o = flag_z[2];
  /* TG68K_ALU.vhd:1042:87  */
  assign n12253_o = {n12251_o, n12252_o};
  /* TG68K_ALU.vhd:1042:97  */
  assign n12255_o = {n12253_o, 2'b00};
  /* TG68K_ALU.vhd:1039:49  */
  assign n12256_o = n12245_o ? n12250_o : n12255_o;
  /* TG68K_ALU.vhd:1037:49  */
  assign n12257_o = v_flag ? 4'b1010 : n12256_o;
  /* TG68K_ALU.vhd:1044:51  */
  assign n12258_o = exec[68];
  /* TG68K_ALU.vhd:1044:72  */
  assign n12260_o = 1'b1 & n12258_o;
  /* TG68K_ALU.vhd:1045:70  */
  assign n12261_o = set_flags[3];
  /* TG68K_ALU.vhd:1046:70  */
  assign n12262_o = set_flags[2];
  /* TG68K_ALU.vhd:1046:83  */
  assign n12263_o = n12821_q[2];
  /* TG68K_ALU.vhd:1046:74  */
  assign n12264_o = n12262_o & n12263_o;
  /* TG68K_ALU.vhd:1049:51  */
  assign n12267_o = exec[67];
  /* TG68K_ALU.vhd:1049:71  */
  assign n12269_o = 1'b1 & n12267_o;
  /* TG68K_ALU.vhd:1050:70  */
  assign n12270_o = set_flags[3];
  /* TG68K_ALU.vhd:1051:70  */
  assign n12271_o = set_flags[2];
  /* TG68K_ALU.vhd:1054:51  */
  assign n12273_o = exec[5];
  /* TG68K_ALU.vhd:1054:70  */
  assign n12274_o = exec[6];
  /* TG68K_ALU.vhd:1054:63  */
  assign n12275_o = n12273_o | n12274_o;
  /* TG68K_ALU.vhd:1054:90  */
  assign n12276_o = exec[7];
  /* TG68K_ALU.vhd:1054:83  */
  assign n12277_o = n12275_o | n12276_o;
  /* TG68K_ALU.vhd:1054:110  */
  assign n12278_o = exec[0];
  /* TG68K_ALU.vhd:1054:103  */
  assign n12279_o = n12277_o | n12278_o;
  /* TG68K_ALU.vhd:1054:131  */
  assign n12280_o = exec[1];
  /* TG68K_ALU.vhd:1054:124  */
  assign n12281_o = n12279_o | n12280_o;
  /* TG68K_ALU.vhd:1054:153  */
  assign n12282_o = exec[15];
  /* TG68K_ALU.vhd:1054:146  */
  assign n12283_o = n12281_o | n12282_o;
  /* TG68K_ALU.vhd:1054:174  */
  assign n12284_o = exec[75];
  /* TG68K_ALU.vhd:1054:167  */
  assign n12285_o = n12283_o | n12284_o;
  /* TG68K_ALU.vhd:1054:194  */
  assign n12286_o = exec[20];
  /* TG68K_ALU.vhd:1054:208  */
  assign n12288_o = 1'b1 & n12286_o;
  /* TG68K_ALU.vhd:1054:186  */
  assign n12289_o = n12285_o | n12288_o;
  /* TG68K_ALU.vhd:1057:56  */
  assign n12292_o = exec[75];
  assign n12293_o = set_flags[3];
  /* TG68K_ALU.vhd:1057:49  */
  assign n12294_o = n12292_o ? bf_nflag : n12293_o;
  assign n12295_o = set_flags[2];
  /* TG68K_ALU.vhd:1060:51  */
  assign n12296_o = exec[9];
  /* TG68K_ALU.vhd:1061:79  */
  assign n12297_o = set_flags[3:2];
  /* TG68K_ALU.vhd:1063:60  */
  assign n12299_o = rot_bits == 2'b00;
  /* TG68K_ALU.vhd:1063:81  */
  assign n12300_o = set_flags[3];
  /* TG68K_ALU.vhd:1063:85  */
  assign n12301_o = n12300_o ^ rot_rot;
  /* TG68K_ALU.vhd:1063:98  */
  assign n12302_o = n12301_o | asl_vflag;
  /* TG68K_ALU.vhd:1063:66  */
  assign n12303_o = n12302_o & n12299_o;
  /* TG68K_ALU.vhd:1063:49  */
  assign n12306_o = n12303_o ? 1'b1 : 1'b0;
  /* TG68K_ALU.vhd:1068:51  */
  assign n12307_o = exec[81];
  /* TG68K_ALU.vhd:1069:79  */
  assign n12308_o = set_flags[3:2];
  /* TG68K_ALU.vhd:1072:51  */
  assign n12309_o = exec[14];
  /* TG68K_ALU.vhd:1073:61  */
  assign n12310_o = ~one_bit_in;
  /* TG68K_ALU.vhd:1074:51  */
  assign n12311_o = exec[87];
  /* TG68K_ALU.vhd:1079:63  */
  assign n12312_o = last_flags1[0];
  /* TG68K_ALU.vhd:1079:66  */
  assign n12313_o = ~n12312_o;
  /* TG68K_ALU.vhd:1080:74  */
  assign n12314_o = n12821_q[0];
  /* TG68K_ALU.vhd:1080:95  */
  assign n12315_o = set_flags[0];
  /* TG68K_ALU.vhd:1080:82  */
  assign n12316_o = ~n12315_o;
  /* TG68K_ALU.vhd:1080:116  */
  assign n12317_o = set_flags[2];
  /* TG68K_ALU.vhd:1080:103  */
  assign n12318_o = ~n12317_o;
  /* TG68K_ALU.vhd:1080:99  */
  assign n12319_o = n12316_o & n12318_o;
  /* TG68K_ALU.vhd:1080:78  */
  assign n12320_o = n12314_o | n12319_o;
  /* TG68K_ALU.vhd:1082:75  */
  assign n12321_o = n12821_q[0];
  /* TG68K_ALU.vhd:1082:92  */
  assign n12322_o = set_flags[0];
  /* TG68K_ALU.vhd:1082:79  */
  assign n12323_o = n12321_o ^ n12322_o;
  /* TG68K_ALU.vhd:1082:111  */
  assign n12324_o = n12821_q[2];
  /* TG68K_ALU.vhd:1082:102  */
  assign n12325_o = ~n12324_o;
  /* TG68K_ALU.vhd:1082:97  */
  assign n12326_o = n12323_o & n12325_o;
  /* TG68K_ALU.vhd:1082:132  */
  assign n12327_o = set_flags[2];
  /* TG68K_ALU.vhd:1082:119  */
  assign n12328_o = ~n12327_o;
  /* TG68K_ALU.vhd:1082:115  */
  assign n12329_o = n12326_o & n12328_o;
  /* TG68K_ALU.vhd:1079:49  */
  assign n12330_o = n12313_o ? n12320_o : n12329_o;
  /* TG68K_ALU.vhd:1085:66  */
  assign n12332_o = n12821_q[2];
  /* TG68K_ALU.vhd:1085:82  */
  assign n12333_o = set_flags[2];
  /* TG68K_ALU.vhd:1085:70  */
  assign n12334_o = n12332_o | n12333_o;
  /* TG68K_ALU.vhd:1086:76  */
  assign n12335_o = last_flags1[0];
  /* TG68K_ALU.vhd:1086:61  */
  assign n12336_o = ~n12335_o;
  /* TG68K_ALU.vhd:1087:51  */
  assign n12337_o = exec[31];
  /* TG68K_ALU.vhd:1088:64  */
  assign n12339_o = exe_datatype == 2'b01;
  /* TG68K_ALU.vhd:1089:75  */
  assign n12340_o = op1out[15];
  /* TG68K_ALU.vhd:1091:75  */
  assign n12341_o = op1out[31];
  /* TG68K_ALU.vhd:1088:49  */
  assign n12342_o = n12339_o ? n12340_o : n12341_o;
  /* TG68K_ALU.vhd:1093:58  */
  assign n12343_o = op1out[15:0];
  /* TG68K_ALU.vhd:1093:71  */
  assign n12345_o = n12343_o == 16'b0000000000000000;
  /* TG68K_ALU.vhd:1093:97  */
  assign n12347_o = exe_datatype == 2'b01;
  /* TG68K_ALU.vhd:1093:112  */
  assign n12348_o = op1out[31:16];
  /* TG68K_ALU.vhd:1093:126  */
  assign n12350_o = n12348_o == 16'b0000000000000000;
  /* TG68K_ALU.vhd:1093:103  */
  assign n12351_o = n12347_o | n12350_o;
  /* TG68K_ALU.vhd:1093:80  */
  assign n12352_o = n12351_o & n12345_o;
  /* TG68K_ALU.vhd:1093:49  */
  assign n12355_o = n12352_o ? 1'b1 : 1'b0;
  assign n12358_o = {n12342_o, n12355_o, 1'b0, 1'b0};
  assign n12359_o = data_read[3:0];
  assign n12360_o = data_read[3:0];
  assign n12361_o = n12821_q[3:0];
  /* TG68K_ALU.vhd:1000:33  */
  assign n12362_o = n12182_o ? n12360_o : n12361_o;
  /* TG68K_ALU.vhd:1003:33  */
  assign n12363_o = n12185_o ? n12359_o : n12362_o;
  /* TG68K_ALU.vhd:1087:41  */
  assign n12364_o = n12337_o ? n12358_o : n12363_o;
  assign n12365_o = {n12336_o, n12334_o, 1'b0, n12330_o};
  /* TG68K_ALU.vhd:1074:41  */
  assign n12366_o = n12311_o ? n12365_o : n12364_o;
  assign n12367_o = n12366_o[1:0];
  assign n12368_o = data_read[1:0];
  assign n12369_o = data_read[1:0];
  assign n12370_o = n12821_q[1:0];
  /* TG68K_ALU.vhd:1000:33  */
  assign n12371_o = n12182_o ? n12369_o : n12370_o;
  /* TG68K_ALU.vhd:1003:33  */
  assign n12372_o = n12185_o ? n12368_o : n12371_o;
  /* TG68K_ALU.vhd:1072:41  */
  assign n12373_o = n12309_o ? n12372_o : n12367_o;
  assign n12374_o = n12366_o[2];
  /* TG68K_ALU.vhd:1072:41  */
  assign n12375_o = n12309_o ? n12310_o : n12374_o;
  assign n12376_o = n12366_o[3];
  assign n12377_o = data_read[3];
  assign n12378_o = data_read[3];
  assign n12379_o = n12821_q[3];
  /* TG68K_ALU.vhd:1000:33  */
  assign n12380_o = n12182_o ? n12378_o : n12379_o;
  /* TG68K_ALU.vhd:1003:33  */
  assign n12381_o = n12185_o ? n12377_o : n12380_o;
  /* TG68K_ALU.vhd:1072:41  */
  assign n12382_o = n12309_o ? n12381_o : n12376_o;
  assign n12383_o = {n12382_o, n12375_o, n12373_o};
  assign n12384_o = {n12308_o, bs_v, bs_c};
  /* TG68K_ALU.vhd:1068:41  */
  assign n12385_o = n12307_o ? n12384_o : n12383_o;
  assign n12386_o = {n12297_o, n12306_o, rot_c};
  /* TG68K_ALU.vhd:1060:41  */
  assign n12387_o = n12296_o ? n12386_o : n12385_o;
  assign n12388_o = {n12294_o, n12295_o, 2'b00};
  /* TG68K_ALU.vhd:1054:41  */
  assign n12389_o = n12289_o ? n12388_o : n12387_o;
  assign n12390_o = {n12270_o, n12271_o, set_mv_flag, 1'b0};
  /* TG68K_ALU.vhd:1049:41  */
  assign n12391_o = n12269_o ? n12390_o : n12389_o;
  assign n12392_o = {n12261_o, n12264_o, 1'b0, 1'b0};
  /* TG68K_ALU.vhd:1044:41  */
  assign n12393_o = n12260_o ? n12392_o : n12391_o;
  /* TG68K_ALU.vhd:1036:41  */
  assign n12394_o = n12241_o ? n12257_o : n12393_o;
  /* TG68K_ALU.vhd:1034:41  */
  assign n12395_o = n12238_o ? set_flags : n12394_o;
  assign n12396_o = {n12235_o, n12395_o};
  assign n12397_o = data_read[4:0];
  assign n12398_o = data_read[4:0];
  assign n12399_o = n12821_q[4:0];
  /* TG68K_ALU.vhd:1000:33  */
  assign n12400_o = n12182_o ? n12398_o : n12399_o;
  /* TG68K_ALU.vhd:1003:33  */
  assign n12401_o = n12185_o ? n12397_o : n12400_o;
  /* TG68K_ALU.vhd:1024:33  */
  assign n12402_o = n12216_o ? n12396_o : n12401_o;
  /* TG68K_ALU.vhd:1024:33  */
  assign n12403_o = n12216_o ? n12217_o : last_flags1;
  assign n12404_o = n12402_o[3:0];
  /* TG68K_ALU.vhd:1014:33  */
  assign n12405_o = z_error ? n12214_o : n12404_o;
  assign n12406_o = n12402_o[4];
  assign n12407_o = data_read[4];
  assign n12408_o = data_read[4];
  assign n12409_o = n12821_q[4];
  /* TG68K_ALU.vhd:1000:33  */
  assign n12410_o = n12182_o ? n12408_o : n12409_o;
  /* TG68K_ALU.vhd:1003:33  */
  assign n12411_o = n12185_o ? n12407_o : n12410_o;
  /* TG68K_ALU.vhd:1014:33  */
  assign n12412_o = z_error ? n12411_o : n12406_o;
  /* TG68K_ALU.vhd:1014:33  */
  assign n12413_o = z_error ? last_flags1 : n12403_o;
  assign n12414_o = {n12412_o, n12405_o};
  assign n12415_o = ccrin[4:0];
  /* TG68K_ALU.vhd:1012:33  */
  assign n12416_o = n12196_o ? n12415_o : n12414_o;
  assign n12417_o = ccrin[7:5];
  assign n12418_o = data_read[7:5];
  assign n12419_o = data_read[7:5];
  assign n12420_o = n12821_q[7:5];
  /* TG68K_ALU.vhd:1000:33  */
  assign n12421_o = n12182_o ? n12419_o : n12420_o;
  /* TG68K_ALU.vhd:1003:33  */
  assign n12422_o = n12185_o ? n12418_o : n12421_o;
  /* TG68K_ALU.vhd:1012:33  */
  assign n12423_o = n12196_o ? n12417_o : n12422_o;
  /* TG68K_ALU.vhd:1012:33  */
  assign n12429_o = n12196_o ? last_flags1 : n12413_o;
  assign n12430_o = {n12423_o, n12416_o};
  /* TG68K_ALU.vhd:999:25  */
  assign n12432_o = clkena_lw ? n12429_o : last_flags1;
  /* TG68K_ALU.vhd:999:25  */
  assign n12433_o = clkena_lw ? n12195_o : asl_vflag;
  /* TG68K_ALU.vhd:997:25  */
  assign n12436_o = reset ? last_flags1 : n12432_o;
  /* TG68K_ALU.vhd:997:25  */
  assign n12437_o = reset ? asl_vflag : n12433_o;
  assign n12439_o = n12434_o[4:0];
  assign n12440_o = n12430_o[4:0];
  assign n12441_o = n12821_q[4:0];
  /* TG68K_ALU.vhd:999:25  */
  assign n12442_o = clkena_lw ? n12440_o : n12441_o;
  /* TG68K_ALU.vhd:997:25  */
  assign n12443_o = reset ? n12439_o : n12442_o;
  assign n12444_o = {3'b000, n12443_o};
  /* TG68K_ALU.vhd:1162:45  */
  assign n12451_o = faktorb[31];
  /* TG68K_ALU.vhd:1162:34  */
  assign n12452_o = n12451_o & signedop;
  /* TG68K_ALU.vhd:1162:55  */
  assign n12453_o = n12452_o | fasign;
  /* TG68K_ALU.vhd:1163:45  */
  assign n12454_o = mulu_reg[63];
  /* TG68K_ALU.vhd:1162:17  */
  assign n12456_o = n12453_o ? n12454_o : 1'b0;
  /* TG68K_ALU.vhd:1168:44  */
  assign n12457_o = faktorb[31];
  /* TG68K_ALU.vhd:1168:33  */
  assign n12458_o = n12457_o & signedop;
  /* TG68K_ALU.vhd:1168:17  */
  assign n12461_o = n12458_o ? 1'b1 : 1'b0;
  /* TG68K_ALU.vhd:1185:70  */
  assign n12462_o = mulu_reg[63:1];
  /* TG68K_ALU.vhd:1185:61  */
  assign n12463_o = {muls_msb, n12462_o};
  /* TG68K_ALU.vhd:1186:36  */
  assign n12464_o = mulu_reg[0];
  /* TG68K_ALU.vhd:1188:88  */
  assign n12465_o = mulu_reg[63:32];
  /* TG68K_ALU.vhd:1188:79  */
  assign n12466_o = {muls_msb, n12465_o};
  /* TG68K_ALU.vhd:1188:113  */
  assign n12467_o = {mulu_sign, faktorb};
  /* TG68K_ALU.vhd:1188:102  */
  assign n12468_o = n12466_o - n12467_o;
  /* TG68K_ALU.vhd:1190:88  */
  assign n12469_o = mulu_reg[63:32];
  /* TG68K_ALU.vhd:1190:79  */
  assign n12470_o = {muls_msb, n12469_o};
  /* TG68K_ALU.vhd:1190:113  */
  assign n12471_o = {mulu_sign, faktorb};
  /* TG68K_ALU.vhd:1190:102  */
  assign n12472_o = n12470_o + n12471_o;
  /* TG68K_ALU.vhd:1187:33  */
  assign n12473_o = fasign ? n12468_o : n12472_o;
  assign n12474_o = n12463_o[63:31];
  /* TG68K_ALU.vhd:1186:25  */
  assign n12475_o = n12464_o ? n12473_o : n12474_o;
  assign n12476_o = n12463_o[30:0];
  /* TG68K_ALU.vhd:1194:30  */
  assign n12477_o = exe_opcode[15];
  /* TG68K_ALU.vhd:1194:39  */
  assign n12479_o = n12477_o | 1'b0;
  /* TG68K_ALU.vhd:1195:56  */
  assign n12480_o = op2out[15:0];
  assign n12482_o = {n12480_o, 16'b0000000000000000};
  /* TG68K_ALU.vhd:1194:17  */
  assign n12483_o = n12479_o ? n12482_o : op2out;
  /* TG68K_ALU.vhd:1201:32  */
  assign n12484_o = result_mulu[63:32];
  /* TG68K_ALU.vhd:1201:46  */
  assign n12486_o = n12484_o == 32'b00000000000000000000000000000000;
  /* TG68K_ALU.vhd:1201:72  */
  assign n12487_o = ~signedop;
  /* TG68K_ALU.vhd:1201:91  */
  assign n12488_o = result_mulu[31];
  /* TG68K_ALU.vhd:1201:95  */
  assign n12489_o = ~n12488_o;
  /* TG68K_ALU.vhd:1201:77  */
  assign n12490_o = n12487_o | n12489_o;
  /* TG68K_ALU.vhd:1201:59  */
  assign n12491_o = n12490_o & n12486_o;
  /* TG68K_ALU.vhd:1202:37  */
  assign n12492_o = result_mulu[63:32];
  /* TG68K_ALU.vhd:1202:51  */
  assign n12494_o = n12492_o == 32'b11111111111111111111111111111111;
  /* TG68K_ALU.vhd:1202:64  */
  assign n12495_o = signedop & n12494_o;
  /* TG68K_ALU.vhd:1202:96  */
  assign n12496_o = result_mulu[31];
  /* TG68K_ALU.vhd:1202:81  */
  assign n12497_o = n12496_o & n12495_o;
  /* TG68K_ALU.vhd:1201:102  */
  assign n12498_o = n12491_o | n12497_o;
  /* TG68K_ALU.vhd:1201:17  */
  assign n12501_o = n12498_o ? 1'b0 : 1'b1;
  /* TG68K_ALU.vhd:1214:55  */
  assign n12507_o = micro_state == 7'b1010101;
  /* TG68K_ALU.vhd:1216:77  */
  assign n12509_o = exe_opcode[15];
  /* TG68K_ALU.vhd:1216:96  */
  assign n12510_o = reg_qa[15];
  /* TG68K_ALU.vhd:1216:86  */
  assign n12511_o = n12510_o & n12509_o;
  /* TG68K_ALU.vhd:1216:120  */
  assign n12512_o = exe_opcode[15];
  /* TG68K_ALU.vhd:1216:124  */
  assign n12513_o = ~n12512_o;
  /* TG68K_ALU.vhd:1216:139  */
  assign n12514_o = reg_qa[31];
  /* TG68K_ALU.vhd:1216:129  */
  assign n12515_o = n12514_o & n12513_o;
  /* TG68K_ALU.vhd:1216:106  */
  assign n12516_o = n12511_o | n12515_o;
  /* TG68K_ALU.vhd:1216:61  */
  assign n12517_o = n12516_o & divs;
  /* TG68K_ALU.vhd:1218:83  */
  assign n12519_o = 32'b00000000000000000000000000000000 - reg_qa;
  /* TG68K_ALU.vhd:1216:49  */
  assign n12520_o = n12517_o ? n12519_o : reg_qa;
  /* TG68K_ALU.vhd:1216:49  */
  assign n12523_o = n12517_o ? 1'b1 : 1'b0;
  /* TG68K_ALU.vhd:1223:51  */
  assign n12524_o = exec[20];
  /* TG68K_ALU.vhd:1223:60  */
  assign n12525_o = ~n12524_o;
  /* TG68K_ALU.vhd:1224:72  */
  assign n12526_o = result_mulu[63:0];
  /* TG68K_ALU.vhd:1223:41  */
  assign n12527_o = n12525_o ? n12526_o : mulu_reg;
  assign n12528_o = {32'b00000000000000000000000000000000, n12520_o};
  /* TG68K_ALU.vhd:1214:41  */
  assign n12529_o = n12507_o ? n12528_o : n12527_o;
  /* TG68K_ALU.vhd:1212:25  */
  assign n12532_o = n12507_o & clkena_lw;
  /* TG68K_ALU.vhd:1240:32  */
  assign n12538_o = opcode[15];
  /* TG68K_ALU.vhd:1240:47  */
  assign n12539_o = opcode[8];
  /* TG68K_ALU.vhd:1240:37  */
  assign n12540_o = n12538_o & n12539_o;
  /* TG68K_ALU.vhd:1240:66  */
  assign n12541_o = opcode[15];
  /* TG68K_ALU.vhd:1240:56  */
  assign n12542_o = ~n12541_o;
  /* TG68K_ALU.vhd:1240:81  */
  assign n12543_o = sndopc[11];
  /* TG68K_ALU.vhd:1240:71  */
  assign n12544_o = n12542_o & n12543_o;
  /* TG68K_ALU.vhd:1240:52  */
  assign n12545_o = n12540_o | n12544_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12547_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12548_o = divs & n12547_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12549_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12550_o = divs & n12549_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12551_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12552_o = divs & n12551_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12553_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12554_o = divs & n12553_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12555_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12556_o = divs & n12555_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12557_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12558_o = divs & n12557_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12559_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12560_o = divs & n12559_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12561_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12562_o = divs & n12561_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12563_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12564_o = divs & n12563_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12565_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12566_o = divs & n12565_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12567_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12568_o = divs & n12567_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12569_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12570_o = divs & n12569_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12571_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12572_o = divs & n12571_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12573_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12574_o = divs & n12573_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12575_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12576_o = divs & n12575_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12577_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12578_o = divs & n12577_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12579_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12580_o = divs & n12579_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12581_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12582_o = divs & n12581_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12583_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12584_o = divs & n12583_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12585_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12586_o = divs & n12585_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12587_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12588_o = divs & n12587_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12589_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12590_o = divs & n12589_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12591_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12592_o = divs & n12591_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12593_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12594_o = divs & n12593_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12595_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12596_o = divs & n12595_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12597_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12598_o = divs & n12597_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12599_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12600_o = divs & n12599_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12601_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12602_o = divs & n12601_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12603_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12604_o = divs & n12603_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12605_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12606_o = divs & n12605_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12607_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12608_o = divs & n12607_o;
  /* TG68K_ALU.vhd:1242:68  */
  assign n12609_o = reg_qa[31];
  /* TG68K_ALU.vhd:1242:58  */
  assign n12610_o = divs & n12609_o;
  assign n12611_o = {n12548_o, n12550_o, n12552_o, n12554_o};
  assign n12612_o = {n12556_o, n12558_o, n12560_o, n12562_o};
  assign n12613_o = {n12564_o, n12566_o, n12568_o, n12570_o};
  assign n12614_o = {n12572_o, n12574_o, n12576_o, n12578_o};
  assign n12615_o = {n12580_o, n12582_o, n12584_o, n12586_o};
  assign n12616_o = {n12588_o, n12590_o, n12592_o, n12594_o};
  assign n12617_o = {n12596_o, n12598_o, n12600_o, n12602_o};
  assign n12618_o = {n12604_o, n12606_o, n12608_o, n12610_o};
  assign n12619_o = {n12611_o, n12612_o, n12613_o, n12614_o};
  assign n12620_o = {n12615_o, n12616_o, n12617_o, n12618_o};
  assign n12621_o = {n12619_o, n12620_o};
  /* TG68K_ALU.vhd:1243:30  */
  assign n12622_o = exe_opcode[15];
  /* TG68K_ALU.vhd:1243:39  */
  assign n12624_o = n12622_o | 1'b0;
  /* TG68K_ALU.vhd:1245:52  */
  assign n12625_o = result_div_pre[15];
  /* TG68K_ALU.vhd:1248:38  */
  assign n12626_o = exe_opcode[14];
  /* TG68K_ALU.vhd:1248:57  */
  assign n12627_o = sndopc[10];
  /* TG68K_ALU.vhd:1248:47  */
  assign n12628_o = n12627_o & n12626_o;
  /* TG68K_ALU.vhd:1248:25  */
  assign n12629_o = n12628_o ? reg_qb : n12621_o;
  /* TG68K_ALU.vhd:1251:52  */
  assign n12630_o = result_div_pre[31];
  /* TG68K_ALU.vhd:1243:17  */
  assign n12631_o = n12624_o ? n12625_o : n12630_o;
  assign n12632_o = {n12629_o, reg_qa};
  assign n12633_o = n12632_o[15:0];
  /* TG68K_ALU.vhd:1243:17  */
  assign n12634_o = n12624_o ? 16'b0000000000000000 : n12633_o;
  assign n12635_o = n12632_o[47:16];
  /* TG68K_ALU.vhd:1243:17  */
  assign n12636_o = n12624_o ? reg_qa : n12635_o;
  assign n12637_o = n12632_o[63:48];
  assign n12638_o = n12621_o[31:16];
  /* TG68K_ALU.vhd:1243:17  */
  assign n12639_o = n12624_o ? n12638_o : n12637_o;
  /* TG68K_ALU.vhd:1253:42  */
  assign n12641_o = opcode[15];
  /* TG68K_ALU.vhd:1253:46  */
  assign n12642_o = ~n12641_o;
  /* TG68K_ALU.vhd:1253:33  */
  assign n12643_o = signedop | n12642_o;
  /* TG68K_ALU.vhd:1254:44  */
  assign n12644_o = op2out[31:16];
  /* TG68K_ALU.vhd:1253:17  */
  assign n12646_o = n12643_o ? n12644_o : 16'b0000000000000000;
  /* TG68K_ALU.vhd:1258:43  */
  assign n12647_o = op2out[31];
  /* TG68K_ALU.vhd:1258:33  */
  assign n12648_o = n12647_o & signedop;
  /* TG68K_ALU.vhd:1259:44  */
  assign n12649_o = div_reg[63:31];
  /* TG68K_ALU.vhd:1259:64  */
  assign n12651_o = {1'b1, op2out};
  /* TG68K_ALU.vhd:1259:59  */
  assign n12652_o = n12649_o + n12651_o;
  /* TG68K_ALU.vhd:1261:44  */
  assign n12653_o = div_reg[63:31];
  /* TG68K_ALU.vhd:1261:64  */
  assign n12655_o = {1'b0, op2outext};
  /* TG68K_ALU.vhd:1261:94  */
  assign n12656_o = op2out[15:0];
  /* TG68K_ALU.vhd:1261:87  */
  assign n12657_o = {n12655_o, n12656_o};
  /* TG68K_ALU.vhd:1261:59  */
  assign n12658_o = n12653_o - n12657_o;
  /* TG68K_ALU.vhd:1258:17  */
  assign n12659_o = n12648_o ? n12652_o : n12658_o;
  /* TG68K_ALU.vhd:1266:43  */
  assign n12660_o = div_sub[32];
  /* TG68K_ALU.vhd:1269:58  */
  assign n12661_o = div_reg[62:31];
  /* TG68K_ALU.vhd:1271:58  */
  assign n12662_o = div_sub[31:0];
  /* TG68K_ALU.vhd:1268:17  */
  assign n12663_o = div_bit ? n12661_o : n12662_o;
  /* TG68K_ALU.vhd:1273:49  */
  assign n12664_o = div_reg[30:0];
  /* TG68K_ALU.vhd:1273:63  */
  assign n12665_o = ~div_bit;
  /* TG68K_ALU.vhd:1273:62  */
  assign n12666_o = {n12664_o, n12665_o};
  /* TG68K_ALU.vhd:1276:66  */
  assign n12667_o = div_quot[31:0];
  /* TG68K_ALU.vhd:1276:57  */
  assign n12669_o = 32'b00000000000000000000000000000000 - n12667_o;
  /* TG68K_ALU.vhd:1279:64  */
  assign n12670_o = div_quot[31:0];
  /* TG68K_ALU.vhd:1275:17  */
  assign n12671_o = div_neg ? n12669_o : n12670_o;
  /* TG68K_ALU.vhd:1282:44  */
  assign n12672_o = ~div_bit;
  /* TG68K_ALU.vhd:1282:34  */
  assign n12673_o = nozero | n12672_o;
  /* TG68K_ALU.vhd:1282:50  */
  assign n12674_o = signedop & n12673_o;
  /* TG68K_ALU.vhd:1282:78  */
  assign n12675_o = op2out[31];
  /* TG68K_ALU.vhd:1282:83  */
  assign n12676_o = n12675_o ^ op1_sign;
  /* TG68K_ALU.vhd:1282:96  */
  assign n12677_o = n12676_o ^ div_qsign;
  /* TG68K_ALU.vhd:1282:67  */
  assign n12678_o = n12677_o & n12674_o;
  /* TG68K_ALU.vhd:1283:37  */
  assign n12679_o = ~signedop;
  /* TG68K_ALU.vhd:1283:54  */
  assign n12680_o = div_over[32];
  /* TG68K_ALU.vhd:1283:58  */
  assign n12681_o = ~n12680_o;
  /* TG68K_ALU.vhd:1283:42  */
  assign n12682_o = n12681_o & n12679_o;
  /* TG68K_ALU.vhd:1283:25  */
  assign n12683_o = n12678_o | n12682_o;
  /* TG68K_ALU.vhd:1283:65  */
  assign n12685_o = 1'b1 & n12683_o;
  /* TG68K_ALU.vhd:1282:17  */
  assign n12688_o = n12685_o ? 1'b1 : 1'b0;
  /* TG68K_ALU.vhd:1294:47  */
  assign n12694_o = micro_state != 7'b1011110;
  /* TG68K_ALU.vhd:1298:47  */
  assign n12697_o = micro_state == 7'b1011001;
  /* TG68K_ALU.vhd:1300:65  */
  assign n12698_o = dividend[63];
  /* TG68K_ALU.vhd:1300:53  */
  assign n12699_o = n12698_o & divs;
  /* TG68K_ALU.vhd:1302:61  */
  assign n12701_o = 64'b0000000000000000000000000000000000000000000000000000000000000000 - dividend;
  /* TG68K_ALU.vhd:1300:41  */
  assign n12702_o = n12699_o ? n12701_o : dividend;
  /* TG68K_ALU.vhd:1300:41  */
  assign n12705_o = n12699_o ? 1'b1 : 1'b0;
  /* TG68K_ALU.vhd:1309:51  */
  assign n12706_o = ~div_bit;
  /* TG68K_ALU.vhd:1309:63  */
  assign n12707_o = n12706_o | nozero;
  /* TG68K_ALU.vhd:1298:33  */
  assign n12708_o = n12697_o ? n12702_o : div_quot;
  /* TG68K_ALU.vhd:1298:33  */
  assign n12710_o = n12697_o ? 1'b0 : n12707_o;
  /* TG68K_ALU.vhd:1311:47  */
  assign n12713_o = micro_state == 7'b1011010;
  /* TG68K_ALU.vhd:1312:72  */
  assign n12714_o = op2out[31];
  /* TG68K_ALU.vhd:1312:77  */
  assign n12715_o = n12714_o ^ op1_sign;
  /* TG68K_ALU.vhd:1312:61  */
  assign n12716_o = signedop & n12715_o;
  /* TG68K_ALU.vhd:1316:73  */
  assign n12717_o = div_reg[63:32];
  /* TG68K_ALU.vhd:1316:65  */
  assign n12719_o = {1'b0, n12717_o};
  /* TG68K_ALU.vhd:1316:93  */
  assign n12721_o = {1'b0, op2outext};
  /* TG68K_ALU.vhd:1316:123  */
  assign n12722_o = op2out[15:0];
  /* TG68K_ALU.vhd:1316:116  */
  assign n12723_o = {n12721_o, n12722_o};
  /* TG68K_ALU.vhd:1316:88  */
  assign n12724_o = n12719_o - n12723_o;
  /* TG68K_ALU.vhd:1319:40  */
  assign n12727_o = exec[68];
  /* TG68K_ALU.vhd:1319:56  */
  assign n12728_o = ~n12727_o;
  /* TG68K_ALU.vhd:1322:87  */
  assign n12729_o = div_quot[63:32];
  /* TG68K_ALU.vhd:1322:78  */
  assign n12731_o = 32'b00000000000000000000000000000000 - n12729_o;
  /* TG68K_ALU.vhd:1324:85  */
  assign n12732_o = div_quot[63:32];
  /* TG68K_ALU.vhd:1321:41  */
  assign n12733_o = op1_sign ? n12731_o : n12732_o;
  assign n12734_o = {n12733_o, result_div_pre};
  /* TG68K_ALU.vhd:1293:25  */
  assign n12736_o = n12728_o & clkena_lw;
  /* TG68K_ALU.vhd:1293:25  */
  assign n12737_o = n12694_o & clkena_lw;
  /* TG68K_ALU.vhd:1293:25  */
  assign n12739_o = n12713_o & clkena_lw;
  /* TG68K_ALU.vhd:1293:25  */
  assign n12740_o = n12713_o & clkena_lw;
  /* TG68K_ALU.vhd:1293:25  */
  assign n12743_o = n12697_o & clkena_lw;
  assign n12753_o = {n9894_o, n9891_o};
  assign n12754_o = {n10045_o, n10038_o, n10031_o};
  assign n12755_o = {n10023_o, n10022_o, n10017_o, n9975_o};
  /* TG68K_ALU.vhd:996:17  */
  always @(posedge clk)
    n12756_q <= n12436_o;
  /* TG68K_ALU.vhd:996:17  */
  assign n12757_o = {n10067_o, n10105_o};
  assign n12759_o = {64'bZ, n12475_o, n12476_o};
  /* TG68K_ALU.vhd:1292:17  */
  assign n12760_o = n12736_o ? n12734_o : result_div;
  /* TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n12761_q <= n12760_o;
  /* TG68K_ALU.vhd:1292:17  */
  assign n12762_o = n12737_o ? n12688_o : v_flag;
  /* TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n12763_q <= n12762_o;
  /* TG68K_ALU.vhd:996:17  */
  always @(posedge clk)
    n12764_q <= n12437_o;
  /* TG68K_ALU.vhd:405:17  */
  assign n12766_o = clkena_lw ? n10126_o : bchg;
  /* TG68K_ALU.vhd:405:17  */
  always @(posedge clk)
    n12767_q <= n12766_o;
  /* TG68K_ALU.vhd:405:17  */
  assign n12768_o = clkena_lw ? n10130_o : bset;
  /* TG68K_ALU.vhd:405:17  */
  always @(posedge clk)
    n12769_q <= n12768_o;
  /* TG68K_ALU.vhd:1211:17  */
  assign n12771_o = clkena_lw ? n12529_o : mulu_reg;
  /* TG68K_ALU.vhd:1211:17  */
  always @(posedge clk)
    n12772_q <= n12771_o;
  /* TG68K_ALU.vhd:1211:17  */
  assign n12773_o = n12532_o ? n12523_o : fasign;
  /* TG68K_ALU.vhd:1211:17  */
  always @(posedge clk)
    n12774_q <= n12773_o;
  /* TG68K_ALU.vhd:1292:17  */
  assign n12776_o = clkena_lw ? n12708_o : div_reg;
  /* TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n12777_q <= n12776_o;
  /* TG68K_ALU.vhd:1292:17  */
  assign n12778_o = {n12663_o, n12666_o};
  /* TG68K_ALU.vhd:1292:17  */
  assign n12780_o = n12739_o ? n12716_o : div_neg;
  /* TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n12781_q <= n12780_o;
  /* TG68K_ALU.vhd:1292:17  */
  assign n12782_o = n12740_o ? n12724_o : div_over;
  /* TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n12783_q <= n12782_o;
  /* TG68K_ALU.vhd:1292:17  */
  assign n12784_o = clkena_lw ? n12710_o : nozero;
  /* TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n12785_q <= n12784_o;
  /* TG68K_ALU.vhd:1292:17  */
  assign n12786_o = {n12639_o, n12636_o, n12634_o};
  /* TG68K_ALU.vhd:1292:17  */
  assign n12787_o = clkena_lw ? divs : signedop;
  /* TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n12788_q <= n12787_o;
  /* TG68K_ALU.vhd:1292:17  */
  assign n12789_o = n12743_o ? n12705_o : op1_sign;
  /* TG68K_ALU.vhd:1292:17  */
  always @(posedge clk)
    n12790_q <= n12789_o;
  assign n12793_o = {n10705_o, n10693_o, n10678_o, n10663_o, n10648_o, n10633_o, n10618_o, n10603_o, n10588_o, n10573_o, n10558_o, n10543_o, n10528_o, n10513_o, n10498_o, n10483_o, n10468_o, n10453_o, n10438_o, n10423_o, n10408_o, n10393_o, n10378_o, n10363_o, n10348_o, n10333_o, n10318_o, n10303_o, n10288_o, n10273_o, n10258_o, n10242_o};
  assign n12795_o = {n11468_o, n11458_o, n11441_o, n11424_o, n11407_o, n11390_o, n11373_o, n11356_o, n11339_o, n11322_o, n11305_o, n11288_o, n11271_o, n11254_o, n11237_o, n11220_o, n11203_o, n11186_o, n11169_o, n11152_o, n11135_o, n11118_o, n11101_o, n11084_o, n11067_o, n11050_o, n11033_o, n11016_o, n10999_o, n10982_o, n10965_o, n10948_o, n10931_o, n10914_o, n10897_o, n10880_o, n10863_o, n10846_o, n10829_o, n10812_o};
  assign n12796_o = {n10706_o, n10698_o, n10683_o, n10668_o, n10653_o, n10638_o, n10623_o, n10608_o, n10593_o, n10578_o, n10563_o, n10548_o, n10533_o, n10518_o, n10503_o, n10488_o, n10473_o, n10458_o, n10443_o, n10428_o, n10413_o, n10398_o, n10383_o, n10368_o, n10353_o, n10338_o, n10323_o, n10308_o, n10293_o, n10278_o, n10263_o, n10247_o};
  assign n12798_o = {n10762_o, n10763_o};
  assign n12799_o = {n11552_o, n11581_o, n11578_o};
  /* TG68K_ALU.vhd:446:17  */
  assign n12800_o = clkena_lw ? n10189_o : bf_bset;
  /* TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n12801_q <= n12800_o;
  /* TG68K_ALU.vhd:446:17  */
  assign n12802_o = clkena_lw ? n10193_o : bf_bchg;
  /* TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n12803_q <= n12802_o;
  /* TG68K_ALU.vhd:446:17  */
  assign n12804_o = clkena_lw ? n10197_o : bf_ins;
  /* TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n12805_q <= n12804_o;
  /* TG68K_ALU.vhd:446:17  */
  assign n12806_o = clkena_lw ? n10201_o : bf_exts;
  /* TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n12807_q <= n12806_o;
  /* TG68K_ALU.vhd:446:17  */
  assign n12808_o = clkena_lw ? n10205_o : bf_fffo;
  /* TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n12809_q <= n12808_o;
  /* TG68K_ALU.vhd:446:17  */
  assign n12810_o = clkena_lw ? n10214_o : bf_d32;
  /* TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n12811_q <= n12810_o;
  /* TG68K_ALU.vhd:446:17  */
  assign n12812_o = clkena_lw ? n10208_o : bf_s32;
  /* TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n12813_q <= n12812_o;
  assign n12815_o = {n12072_o, n12070_o, n12067_o, n12064_o, n12061_o, n12074_o};
  assign n12816_o = {n11753_o, n11750_o, n11754_o, n11748_o, n11752_o};
  assign n12817_o = {n12007_o, n12009_o};
  assign n12818_o = {n12088_o, n12083_o, n12094_o};
  /* TG68K_ALU.vhd:446:17  */
  assign n12819_o = clkena_lw ? n10216_o : n12820_q;
  /* TG68K_ALU.vhd:446:17  */
  always @(posedge clk)
    n12820_q <= n12819_o;
  /* TG68K_ALU.vhd:996:17  */
  always @(posedge clk)
    n12821_q <= n12444_o;
  /* TG68K_ALU.vhd:76:17  */
  assign n12822_o = op1out[0];
  /* TG68K_ALU.vhd:75:17  */
  assign n12823_o = op1out[1];
  /* TG68K_ALU.vhd:74:17  */
  assign n12824_o = op1out[2];
  /* TG68K_ALU.vhd:73:17  */
  assign n12825_o = op1out[3];
  /* TG68K_ALU.vhd:72:17  */
  assign n12826_o = op1out[4];
  /* TG68K_ALU.vhd:66:17  */
  assign n12827_o = op1out[5];
  /* TG68K_ALU.vhd:446:17  */
  assign n12828_o = op1out[6];
  assign n12829_o = op1out[7];
  assign n12830_o = op1out[8];
  assign n12831_o = op1out[9];
  /* TG68K_ALU.vhd:1292:17  */
  assign n12832_o = op1out[10];
  assign n12833_o = op1out[11];
  /* TG68K_ALU.vhd:1211:17  */
  assign n12834_o = op1out[12];
  /* TG68K_ALU.vhd:405:17  */
  assign n12835_o = op1out[13];
  /* TG68K_ALU.vhd:996:17  */
  assign n12836_o = op1out[14];
  assign n12837_o = op1out[15];
  /* TG68K_ALU.vhd:1292:17  */
  assign n12838_o = op1out[16];
  /* TG68K_ALU.vhd:1292:17  */
  assign n12839_o = op1out[17];
  /* TG68K_ALU.vhd:1292:17  */
  assign n12840_o = op1out[18];
  /* TG68K_ALU.vhd:1292:17  */
  assign n12841_o = op1out[19];
  /* TG68K_ALU.vhd:1292:17  */
  assign n12842_o = op1out[20];
  /* TG68K_ALU.vhd:1292:17  */
  assign n12843_o = op1out[21];
  /* TG68K_ALU.vhd:1292:17  */
  assign n12844_o = op1out[22];
  /* TG68K_ALU.vhd:1292:17  */
  assign n12845_o = op1out[23];
  /* TG68K_ALU.vhd:1290:1  */
  assign n12846_o = op1out[24];
  assign n12847_o = op1out[25];
  assign n12848_o = op1out[26];
  /* TG68K_ALU.vhd:1237:1  */
  assign n12849_o = op1out[27];
  assign n12850_o = op1out[28];
  /* TG68K_ALU.vhd:1211:17  */
  assign n12851_o = op1out[29];
  /* TG68K_ALU.vhd:1211:17  */
  assign n12852_o = op1out[30];
  /* TG68K_ALU.vhd:1209:1  */
  assign n12853_o = op1out[31];
  /* TG68K_ALU.vhd:433:37  */
  assign n12854_o = bit_number[1:0];
  /* TG68K_ALU.vhd:433:37  */
  always @*
    case (n12854_o)
      2'b00: n12855_o = n12822_o;
      2'b01: n12855_o = n12823_o;
      2'b10: n12855_o = n12824_o;
      2'b11: n12855_o = n12825_o;
    endcase
  /* TG68K_ALU.vhd:433:37  */
  assign n12856_o = bit_number[1:0];
  /* TG68K_ALU.vhd:433:37  */
  always @*
    case (n12856_o)
      2'b00: n12857_o = n12826_o;
      2'b01: n12857_o = n12827_o;
      2'b10: n12857_o = n12828_o;
      2'b11: n12857_o = n12829_o;
    endcase
  /* TG68K_ALU.vhd:433:37  */
  assign n12858_o = bit_number[1:0];
  /* TG68K_ALU.vhd:433:37  */
  always @*
    case (n12858_o)
      2'b00: n12859_o = n12830_o;
      2'b01: n12859_o = n12831_o;
      2'b10: n12859_o = n12832_o;
      2'b11: n12859_o = n12833_o;
    endcase
  /* TG68K_ALU.vhd:433:37  */
  assign n12860_o = bit_number[1:0];
  /* TG68K_ALU.vhd:433:37  */
  always @*
    case (n12860_o)
      2'b00: n12861_o = n12834_o;
      2'b01: n12861_o = n12835_o;
      2'b10: n12861_o = n12836_o;
      2'b11: n12861_o = n12837_o;
    endcase
  /* TG68K_ALU.vhd:433:37  */
  assign n12862_o = bit_number[1:0];
  /* TG68K_ALU.vhd:433:37  */
  always @*
    case (n12862_o)
      2'b00: n12863_o = n12838_o;
      2'b01: n12863_o = n12839_o;
      2'b10: n12863_o = n12840_o;
      2'b11: n12863_o = n12841_o;
    endcase
  /* TG68K_ALU.vhd:433:37  */
  assign n12864_o = bit_number[1:0];
  /* TG68K_ALU.vhd:433:37  */
  always @*
    case (n12864_o)
      2'b00: n12865_o = n12842_o;
      2'b01: n12865_o = n12843_o;
      2'b10: n12865_o = n12844_o;
      2'b11: n12865_o = n12845_o;
    endcase
  /* TG68K_ALU.vhd:433:37  */
  assign n12866_o = bit_number[1:0];
  /* TG68K_ALU.vhd:433:37  */
  always @*
    case (n12866_o)
      2'b00: n12867_o = n12846_o;
      2'b01: n12867_o = n12847_o;
      2'b10: n12867_o = n12848_o;
      2'b11: n12867_o = n12849_o;
    endcase
  /* TG68K_ALU.vhd:433:37  */
  assign n12868_o = bit_number[1:0];
  /* TG68K_ALU.vhd:433:37  */
  always @*
    case (n12868_o)
      2'b00: n12869_o = n12850_o;
      2'b01: n12869_o = n12851_o;
      2'b10: n12869_o = n12852_o;
      2'b11: n12869_o = n12853_o;
    endcase
  /* TG68K_ALU.vhd:433:37  */
  assign n12870_o = bit_number[3:2];
  /* TG68K_ALU.vhd:433:37  */
  always @*
    case (n12870_o)
      2'b00: n12871_o = n12855_o;
      2'b01: n12871_o = n12857_o;
      2'b10: n12871_o = n12859_o;
      2'b11: n12871_o = n12861_o;
    endcase
  /* TG68K_ALU.vhd:433:37  */
  assign n12872_o = bit_number[3:2];
  /* TG68K_ALU.vhd:433:37  */
  always @*
    case (n12872_o)
      2'b00: n12873_o = n12863_o;
      2'b01: n12873_o = n12865_o;
      2'b10: n12873_o = n12867_o;
      2'b11: n12873_o = n12869_o;
    endcase
  /* TG68K_ALU.vhd:433:37  */
  assign n12874_o = bit_number[4];
  /* TG68K_ALU.vhd:433:37  */
  assign n12875_o = n12874_o ? n12873_o : n12871_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12876_o = bit_number[4];
  /* TG68K_ALU.vhd:435:17  */
  assign n12877_o = ~n12876_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12878_o = bit_number[3];
  /* TG68K_ALU.vhd:435:17  */
  assign n12879_o = ~n12878_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12880_o = n12877_o & n12879_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12881_o = n12877_o & n12878_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12882_o = n12876_o & n12879_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12883_o = n12876_o & n12878_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12884_o = bit_number[2];
  /* TG68K_ALU.vhd:435:17  */
  assign n12885_o = ~n12884_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12886_o = n12880_o & n12885_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12887_o = n12880_o & n12884_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12888_o = n12881_o & n12885_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12889_o = n12881_o & n12884_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12890_o = n12882_o & n12885_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12891_o = n12882_o & n12884_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12892_o = n12883_o & n12885_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12893_o = n12883_o & n12884_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12894_o = bit_number[1];
  /* TG68K_ALU.vhd:435:17  */
  assign n12895_o = ~n12894_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12896_o = n12886_o & n12895_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12897_o = n12886_o & n12894_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12898_o = n12887_o & n12895_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12899_o = n12887_o & n12894_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12900_o = n12888_o & n12895_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12901_o = n12888_o & n12894_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12902_o = n12889_o & n12895_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12903_o = n12889_o & n12894_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12904_o = n12890_o & n12895_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12905_o = n12890_o & n12894_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12906_o = n12891_o & n12895_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12907_o = n12891_o & n12894_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12908_o = n12892_o & n12895_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12909_o = n12892_o & n12894_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12910_o = n12893_o & n12895_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12911_o = n12893_o & n12894_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12912_o = bit_number[0];
  /* TG68K_ALU.vhd:435:17  */
  assign n12913_o = ~n12912_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12914_o = n12896_o & n12913_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12915_o = n12896_o & n12912_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12916_o = n12897_o & n12913_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12917_o = n12897_o & n12912_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12918_o = n12898_o & n12913_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12919_o = n12898_o & n12912_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12920_o = n12899_o & n12913_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12921_o = n12899_o & n12912_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12922_o = n12900_o & n12913_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12923_o = n12900_o & n12912_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12924_o = n12901_o & n12913_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12925_o = n12901_o & n12912_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12926_o = n12902_o & n12913_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12927_o = n12902_o & n12912_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12928_o = n12903_o & n12913_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12929_o = n12903_o & n12912_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12930_o = n12904_o & n12913_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12931_o = n12904_o & n12912_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12932_o = n12905_o & n12913_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12933_o = n12905_o & n12912_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12934_o = n12906_o & n12913_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12935_o = n12906_o & n12912_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12936_o = n12907_o & n12913_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12937_o = n12907_o & n12912_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12938_o = n12908_o & n12913_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12939_o = n12908_o & n12912_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12940_o = n12909_o & n12913_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12941_o = n12909_o & n12912_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12942_o = n12910_o & n12913_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12943_o = n12910_o & n12912_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12944_o = n12911_o & n12913_o;
  /* TG68K_ALU.vhd:435:17  */
  assign n12945_o = n12911_o & n12912_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n12946_o = op1out[0];
  /* TG68K_ALU.vhd:435:17  */
  assign n12947_o = n12914_o ? n10162_o : n12946_o;
  /* TG68K_ALU.vhd:575:17  */
  assign n12948_o = op1out[1];
  /* TG68K_ALU.vhd:435:17  */
  assign n12949_o = n12915_o ? n10162_o : n12948_o;
  assign n12950_o = op1out[2];
  /* TG68K_ALU.vhd:435:17  */
  assign n12951_o = n12916_o ? n10162_o : n12950_o;
  assign n12952_o = op1out[3];
  /* TG68K_ALU.vhd:435:17  */
  assign n12953_o = n12917_o ? n10162_o : n12952_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n12954_o = op1out[4];
  /* TG68K_ALU.vhd:435:17  */
  assign n12955_o = n12918_o ? n10162_o : n12954_o;
  assign n12956_o = op1out[5];
  /* TG68K_ALU.vhd:435:17  */
  assign n12957_o = n12919_o ? n10162_o : n12956_o;
  assign n12958_o = op1out[6];
  /* TG68K_ALU.vhd:435:17  */
  assign n12959_o = n12920_o ? n10162_o : n12958_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n12960_o = op1out[7];
  /* TG68K_ALU.vhd:435:17  */
  assign n12961_o = n12921_o ? n10162_o : n12960_o;
  /* TG68K_ALU.vhd:575:17  */
  assign n12962_o = op1out[8];
  /* TG68K_ALU.vhd:435:17  */
  assign n12963_o = n12922_o ? n10162_o : n12962_o;
  assign n12964_o = op1out[9];
  /* TG68K_ALU.vhd:435:17  */
  assign n12965_o = n12923_o ? n10162_o : n12964_o;
  assign n12966_o = op1out[10];
  /* TG68K_ALU.vhd:435:17  */
  assign n12967_o = n12924_o ? n10162_o : n12966_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n12968_o = op1out[11];
  /* TG68K_ALU.vhd:435:17  */
  assign n12969_o = n12925_o ? n10162_o : n12968_o;
  assign n12970_o = op1out[12];
  /* TG68K_ALU.vhd:435:17  */
  assign n12971_o = n12926_o ? n10162_o : n12970_o;
  assign n12972_o = op1out[13];
  /* TG68K_ALU.vhd:435:17  */
  assign n12973_o = n12927_o ? n10162_o : n12972_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n12974_o = op1out[14];
  /* TG68K_ALU.vhd:435:17  */
  assign n12975_o = n12928_o ? n10162_o : n12974_o;
  /* TG68K_ALU.vhd:575:17  */
  assign n12976_o = op1out[15];
  /* TG68K_ALU.vhd:435:17  */
  assign n12977_o = n12929_o ? n10162_o : n12976_o;
  assign n12978_o = op1out[16];
  /* TG68K_ALU.vhd:435:17  */
  assign n12979_o = n12930_o ? n10162_o : n12978_o;
  assign n12980_o = op1out[17];
  /* TG68K_ALU.vhd:435:17  */
  assign n12981_o = n12931_o ? n10162_o : n12980_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n12982_o = op1out[18];
  /* TG68K_ALU.vhd:435:17  */
  assign n12983_o = n12932_o ? n10162_o : n12982_o;
  assign n12984_o = op1out[19];
  /* TG68K_ALU.vhd:435:17  */
  assign n12985_o = n12933_o ? n10162_o : n12984_o;
  assign n12986_o = op1out[20];
  /* TG68K_ALU.vhd:435:17  */
  assign n12987_o = n12934_o ? n10162_o : n12986_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n12988_o = op1out[21];
  /* TG68K_ALU.vhd:435:17  */
  assign n12989_o = n12935_o ? n10162_o : n12988_o;
  /* TG68K_ALU.vhd:575:17  */
  assign n12990_o = op1out[22];
  /* TG68K_ALU.vhd:435:17  */
  assign n12991_o = n12936_o ? n10162_o : n12990_o;
  assign n12992_o = op1out[23];
  /* TG68K_ALU.vhd:435:17  */
  assign n12993_o = n12937_o ? n10162_o : n12992_o;
  assign n12994_o = op1out[24];
  /* TG68K_ALU.vhd:435:17  */
  assign n12995_o = n12938_o ? n10162_o : n12994_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n12996_o = op1out[25];
  /* TG68K_ALU.vhd:435:17  */
  assign n12997_o = n12939_o ? n10162_o : n12996_o;
  assign n12998_o = op1out[26];
  /* TG68K_ALU.vhd:435:17  */
  assign n12999_o = n12940_o ? n10162_o : n12998_o;
  assign n13000_o = op1out[27];
  /* TG68K_ALU.vhd:435:17  */
  assign n13001_o = n12941_o ? n10162_o : n13000_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n13002_o = op1out[28];
  /* TG68K_ALU.vhd:435:17  */
  assign n13003_o = n12942_o ? n10162_o : n13002_o;
  /* TG68K_ALU.vhd:575:17  */
  assign n13004_o = op1out[29];
  /* TG68K_ALU.vhd:435:17  */
  assign n13005_o = n12943_o ? n10162_o : n13004_o;
  assign n13006_o = op1out[30];
  /* TG68K_ALU.vhd:435:17  */
  assign n13007_o = n12944_o ? n10162_o : n13006_o;
  assign n13008_o = op1out[31];
  /* TG68K_ALU.vhd:435:17  */
  assign n13009_o = n12945_o ? n10162_o : n13008_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n13010_o = {n13009_o, n13007_o, n13005_o, n13003_o, n13001_o, n12999_o, n12997_o, n12995_o, n12993_o, n12991_o, n12989_o, n12987_o, n12985_o, n12983_o, n12981_o, n12979_o, n12977_o, n12975_o, n12973_o, n12971_o, n12969_o, n12967_o, n12965_o, n12963_o, n12961_o, n12959_o, n12957_o, n12955_o, n12953_o, n12951_o, n12949_o, n12947_o};
  /* TG68K_ALU.vhd:435:26  */
  assign n13011_o = datareg[0];
  /* TG68K_ALU.vhd:435:17  */
  assign n13012_o = datareg[1];
  /* TG68K_ALU.vhd:575:17  */
  assign n13013_o = datareg[2];
  assign n13014_o = datareg[3];
  assign n13015_o = datareg[4];
  assign n13016_o = datareg[5];
  assign n13017_o = datareg[6];
  /* TG68K_ALU.vhd:581:17  */
  assign n13018_o = datareg[7];
  /* TG68K_ALU.vhd:572:17  */
  assign n13019_o = datareg[8];
  /* TG68K_ALU.vhd:575:17  */
  assign n13020_o = datareg[9];
  assign n13021_o = datareg[10];
  assign n13022_o = datareg[11];
  assign n13023_o = datareg[12];
  assign n13024_o = datareg[13];
  /* TG68K_ALU.vhd:581:17  */
  assign n13025_o = datareg[14];
  /* TG68K_ALU.vhd:572:17  */
  assign n13026_o = datareg[15];
  /* TG68K_ALU.vhd:575:17  */
  assign n13027_o = datareg[16];
  assign n13028_o = datareg[17];
  assign n13029_o = datareg[18];
  assign n13030_o = datareg[19];
  assign n13031_o = datareg[20];
  /* TG68K_ALU.vhd:581:17  */
  assign n13032_o = datareg[21];
  /* TG68K_ALU.vhd:572:17  */
  assign n13033_o = datareg[22];
  /* TG68K_ALU.vhd:575:17  */
  assign n13034_o = datareg[23];
  assign n13035_o = datareg[24];
  assign n13036_o = datareg[25];
  assign n13037_o = datareg[26];
  assign n13038_o = datareg[27];
  /* TG68K_ALU.vhd:581:17  */
  assign n13039_o = datareg[28];
  /* TG68K_ALU.vhd:572:17  */
  assign n13040_o = datareg[29];
  /* TG68K_ALU.vhd:575:17  */
  assign n13041_o = datareg[30];
  assign n13042_o = datareg[31];
  /* TG68K_ALU.vhd:496:36  */
  assign n13043_o = n10708_o[1:0];
  /* TG68K_ALU.vhd:496:36  */
  always @*
    case (n13043_o)
      2'b00: n13044_o = n13011_o;
      2'b01: n13044_o = n13012_o;
      2'b10: n13044_o = n13013_o;
      2'b11: n13044_o = n13014_o;
    endcase
  /* TG68K_ALU.vhd:496:36  */
  assign n13045_o = n10708_o[1:0];
  /* TG68K_ALU.vhd:496:36  */
  always @*
    case (n13045_o)
      2'b00: n13046_o = n13015_o;
      2'b01: n13046_o = n13016_o;
      2'b10: n13046_o = n13017_o;
      2'b11: n13046_o = n13018_o;
    endcase
  /* TG68K_ALU.vhd:496:36  */
  assign n13047_o = n10708_o[1:0];
  /* TG68K_ALU.vhd:496:36  */
  always @*
    case (n13047_o)
      2'b00: n13048_o = n13019_o;
      2'b01: n13048_o = n13020_o;
      2'b10: n13048_o = n13021_o;
      2'b11: n13048_o = n13022_o;
    endcase
  /* TG68K_ALU.vhd:496:36  */
  assign n13049_o = n10708_o[1:0];
  /* TG68K_ALU.vhd:496:36  */
  always @*
    case (n13049_o)
      2'b00: n13050_o = n13023_o;
      2'b01: n13050_o = n13024_o;
      2'b10: n13050_o = n13025_o;
      2'b11: n13050_o = n13026_o;
    endcase
  /* TG68K_ALU.vhd:496:36  */
  assign n13051_o = n10708_o[1:0];
  /* TG68K_ALU.vhd:496:36  */
  always @*
    case (n13051_o)
      2'b00: n13052_o = n13027_o;
      2'b01: n13052_o = n13028_o;
      2'b10: n13052_o = n13029_o;
      2'b11: n13052_o = n13030_o;
    endcase
  /* TG68K_ALU.vhd:496:36  */
  assign n13053_o = n10708_o[1:0];
  /* TG68K_ALU.vhd:496:36  */
  always @*
    case (n13053_o)
      2'b00: n13054_o = n13031_o;
      2'b01: n13054_o = n13032_o;
      2'b10: n13054_o = n13033_o;
      2'b11: n13054_o = n13034_o;
    endcase
  /* TG68K_ALU.vhd:496:36  */
  assign n13055_o = n10708_o[1:0];
  /* TG68K_ALU.vhd:496:36  */
  always @*
    case (n13055_o)
      2'b00: n13056_o = n13035_o;
      2'b01: n13056_o = n13036_o;
      2'b10: n13056_o = n13037_o;
      2'b11: n13056_o = n13038_o;
    endcase
  /* TG68K_ALU.vhd:496:36  */
  assign n13057_o = n10708_o[1:0];
  /* TG68K_ALU.vhd:496:36  */
  always @*
    case (n13057_o)
      2'b00: n13058_o = n13039_o;
      2'b01: n13058_o = n13040_o;
      2'b10: n13058_o = n13041_o;
      2'b11: n13058_o = n13042_o;
    endcase
  /* TG68K_ALU.vhd:496:36  */
  assign n13059_o = n10708_o[3:2];
  /* TG68K_ALU.vhd:496:36  */
  always @*
    case (n13059_o)
      2'b00: n13060_o = n13044_o;
      2'b01: n13060_o = n13046_o;
      2'b10: n13060_o = n13048_o;
      2'b11: n13060_o = n13050_o;
    endcase
  /* TG68K_ALU.vhd:496:36  */
  assign n13061_o = n10708_o[3:2];
  /* TG68K_ALU.vhd:496:36  */
  always @*
    case (n13061_o)
      2'b00: n13062_o = n13052_o;
      2'b01: n13062_o = n13054_o;
      2'b10: n13062_o = n13056_o;
      2'b11: n13062_o = n13058_o;
    endcase
  /* TG68K_ALU.vhd:496:36  */
  assign n13063_o = n10708_o[4];
  /* TG68K_ALU.vhd:496:36  */
  assign n13064_o = n13063_o ? n13062_o : n13060_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13065_o = bit_msb[5];
  /* TG68K_ALU.vhd:761:17  */
  assign n13066_o = ~n13065_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13067_o = bit_msb[4];
  /* TG68K_ALU.vhd:761:17  */
  assign n13068_o = ~n13067_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13069_o = n13066_o & n13068_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13070_o = n13066_o & n13067_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13071_o = n13065_o & n13068_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13072_o = bit_msb[3];
  /* TG68K_ALU.vhd:761:17  */
  assign n13073_o = ~n13072_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13074_o = n13069_o & n13073_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13075_o = n13069_o & n13072_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13076_o = n13070_o & n13073_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13077_o = n13070_o & n13072_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13078_o = n13071_o & n13073_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13079_o = bit_msb[2];
  /* TG68K_ALU.vhd:761:17  */
  assign n13080_o = ~n13079_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13081_o = n13074_o & n13080_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13082_o = n13074_o & n13079_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13083_o = n13075_o & n13080_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13084_o = n13075_o & n13079_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13085_o = n13076_o & n13080_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13086_o = n13076_o & n13079_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13087_o = n13077_o & n13080_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13088_o = n13077_o & n13079_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13089_o = n13078_o & n13080_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13090_o = bit_msb[1];
  /* TG68K_ALU.vhd:761:17  */
  assign n13091_o = ~n13090_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13092_o = n13081_o & n13091_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13093_o = n13081_o & n13090_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13094_o = n13082_o & n13091_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13095_o = n13082_o & n13090_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13096_o = n13083_o & n13091_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13097_o = n13083_o & n13090_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13098_o = n13084_o & n13091_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13099_o = n13084_o & n13090_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13100_o = n13085_o & n13091_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13101_o = n13085_o & n13090_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13102_o = n13086_o & n13091_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13103_o = n13086_o & n13090_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13104_o = n13087_o & n13091_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13105_o = n13087_o & n13090_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13106_o = n13088_o & n13091_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13107_o = n13088_o & n13090_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13108_o = n13089_o & n13091_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13109_o = bit_msb[0];
  /* TG68K_ALU.vhd:761:17  */
  assign n13110_o = ~n13109_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13111_o = n13092_o & n13110_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13112_o = n13092_o & n13109_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13113_o = n13093_o & n13110_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13114_o = n13093_o & n13109_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13115_o = n13094_o & n13110_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13116_o = n13094_o & n13109_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13117_o = n13095_o & n13110_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13118_o = n13095_o & n13109_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13119_o = n13096_o & n13110_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13120_o = n13096_o & n13109_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13121_o = n13097_o & n13110_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13122_o = n13097_o & n13109_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13123_o = n13098_o & n13110_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13124_o = n13098_o & n13109_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13125_o = n13099_o & n13110_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13126_o = n13099_o & n13109_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13127_o = n13100_o & n13110_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13128_o = n13100_o & n13109_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13129_o = n13101_o & n13110_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13130_o = n13101_o & n13109_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13131_o = n13102_o & n13110_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13132_o = n13102_o & n13109_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13133_o = n13103_o & n13110_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13134_o = n13103_o & n13109_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13135_o = n13104_o & n13110_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13136_o = n13104_o & n13109_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13137_o = n13105_o & n13110_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13138_o = n13105_o & n13109_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13139_o = n13106_o & n13110_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13140_o = n13106_o & n13109_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13141_o = n13107_o & n13110_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13142_o = n13107_o & n13109_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13143_o = n13108_o & n13110_o;
  /* TG68K_ALU.vhd:761:17  */
  assign n13144_o = n13108_o & n13109_o;
  assign n13145_o = n11719_o[0];
  /* TG68K_ALU.vhd:761:17  */
  assign n13146_o = n13111_o ? 1'b1 : n13145_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n13147_o = n11719_o[1];
  /* TG68K_ALU.vhd:761:17  */
  assign n13148_o = n13112_o ? 1'b1 : n13147_o;
  assign n13149_o = n11719_o[2];
  /* TG68K_ALU.vhd:761:17  */
  assign n13150_o = n13113_o ? 1'b1 : n13149_o;
  assign n13151_o = n11719_o[3];
  /* TG68K_ALU.vhd:761:17  */
  assign n13152_o = n13114_o ? 1'b1 : n13151_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n13153_o = n11719_o[4];
  /* TG68K_ALU.vhd:761:17  */
  assign n13154_o = n13115_o ? 1'b1 : n13153_o;
  /* TG68K_ALU.vhd:575:17  */
  assign n13155_o = n11719_o[5];
  /* TG68K_ALU.vhd:761:17  */
  assign n13156_o = n13116_o ? 1'b1 : n13155_o;
  assign n13157_o = n11719_o[6];
  /* TG68K_ALU.vhd:761:17  */
  assign n13158_o = n13117_o ? 1'b1 : n13157_o;
  assign n13159_o = n11719_o[7];
  /* TG68K_ALU.vhd:761:17  */
  assign n13160_o = n13118_o ? 1'b1 : n13159_o;
  /* TG68K_ALU.vhd:572:17  */
  assign n13161_o = n11719_o[8];
  /* TG68K_ALU.vhd:761:17  */
  assign n13162_o = n13119_o ? 1'b1 : n13161_o;
  assign n13163_o = n11719_o[9];
  /* TG68K_ALU.vhd:761:17  */
  assign n13164_o = n13120_o ? 1'b1 : n13163_o;
  assign n13165_o = n11719_o[10];
  /* TG68K_ALU.vhd:761:17  */
  assign n13166_o = n13121_o ? 1'b1 : n13165_o;
  /* TG68K_ALU.vhd:581:17  */
  assign n13167_o = n11719_o[11];
  /* TG68K_ALU.vhd:761:17  */
  assign n13168_o = n13122_o ? 1'b1 : n13167_o;
  /* TG68K_ALU.vhd:575:17  */
  assign n13169_o = n11719_o[12];
  /* TG68K_ALU.vhd:761:17  */
  assign n13170_o = n13123_o ? 1'b1 : n13169_o;
  assign n13171_o = n11719_o[13];
  /* TG68K_ALU.vhd:761:17  */
  assign n13172_o = n13124_o ? 1'b1 : n13171_o;
  assign n13173_o = n11719_o[14];
  /* TG68K_ALU.vhd:761:17  */
  assign n13174_o = n13125_o ? 1'b1 : n13173_o;
  assign n13175_o = n11719_o[15];
  /* TG68K_ALU.vhd:761:17  */
  assign n13176_o = n13126_o ? 1'b1 : n13175_o;
  assign n13177_o = n11719_o[16];
  /* TG68K_ALU.vhd:761:17  */
  assign n13178_o = n13127_o ? 1'b1 : n13177_o;
  assign n13179_o = n11719_o[17];
  /* TG68K_ALU.vhd:761:17  */
  assign n13180_o = n13128_o ? 1'b1 : n13179_o;
  assign n13181_o = n11719_o[18];
  /* TG68K_ALU.vhd:761:17  */
  assign n13182_o = n13129_o ? 1'b1 : n13181_o;
  assign n13183_o = n11719_o[19];
  /* TG68K_ALU.vhd:761:17  */
  assign n13184_o = n13130_o ? 1'b1 : n13183_o;
  assign n13185_o = n11719_o[20];
  /* TG68K_ALU.vhd:761:17  */
  assign n13186_o = n13131_o ? 1'b1 : n13185_o;
  assign n13187_o = n11719_o[21];
  /* TG68K_ALU.vhd:761:17  */
  assign n13188_o = n13132_o ? 1'b1 : n13187_o;
  assign n13189_o = n11719_o[22];
  /* TG68K_ALU.vhd:761:17  */
  assign n13190_o = n13133_o ? 1'b1 : n13189_o;
  assign n13191_o = n11719_o[23];
  /* TG68K_ALU.vhd:761:17  */
  assign n13192_o = n13134_o ? 1'b1 : n13191_o;
  assign n13193_o = n11719_o[24];
  /* TG68K_ALU.vhd:761:17  */
  assign n13194_o = n13135_o ? 1'b1 : n13193_o;
  assign n13195_o = n11719_o[25];
  /* TG68K_ALU.vhd:761:17  */
  assign n13196_o = n13136_o ? 1'b1 : n13195_o;
  assign n13197_o = n11719_o[26];
  /* TG68K_ALU.vhd:761:17  */
  assign n13198_o = n13137_o ? 1'b1 : n13197_o;
  assign n13199_o = n11719_o[27];
  /* TG68K_ALU.vhd:761:17  */
  assign n13200_o = n13138_o ? 1'b1 : n13199_o;
  assign n13201_o = n11719_o[28];
  /* TG68K_ALU.vhd:761:17  */
  assign n13202_o = n13139_o ? 1'b1 : n13201_o;
  assign n13203_o = n11719_o[29];
  /* TG68K_ALU.vhd:761:17  */
  assign n13204_o = n13140_o ? 1'b1 : n13203_o;
  assign n13205_o = n11719_o[30];
  /* TG68K_ALU.vhd:761:17  */
  assign n13206_o = n13141_o ? 1'b1 : n13205_o;
  assign n13207_o = n11719_o[31];
  /* TG68K_ALU.vhd:761:17  */
  assign n13208_o = n13142_o ? 1'b1 : n13207_o;
  assign n13209_o = n11719_o[32];
  /* TG68K_ALU.vhd:761:17  */
  assign n13210_o = n13143_o ? 1'b1 : n13209_o;
  assign n13211_o = n11719_o[33];
  /* TG68K_ALU.vhd:761:17  */
  assign n13212_o = n13144_o ? 1'b1 : n13211_o;
  assign n13213_o = {n13212_o, n13210_o, n13208_o, n13206_o, n13204_o, n13202_o, n13200_o, n13198_o, n13196_o, n13194_o, n13192_o, n13190_o, n13188_o, n13186_o, n13184_o, n13182_o, n13180_o, n13178_o, n13176_o, n13174_o, n13172_o, n13170_o, n13168_o, n13166_o, n13164_o, n13162_o, n13160_o, n13158_o, n13156_o, n13154_o, n13152_o, n13150_o, n13148_o, n13146_o};
endmodule

module tg68kdotc_kernel_0_2_2_2_2_2_0_0
  (input  clk,
   input  nreset,
   input  clkena_in,
   input  [15:0] data_in,
   input  [2:0] ipl,
   input  ipl_autovector,
   input  berr,
   input  [1:0] cpu,
   output [31:0] addr_out,
   output [15:0] data_write,
   output nwr,
   output nuds,
   output nlds,
   output [1:0] busstate,
   output longword,
   output nresetout,
   output [2:0] fc,
   output clr_berr,
   output skipfetch,
   output [31:0] regin_out,
   output [3:0] cacr_out,
   output [31:0] vbr_out);
  wire use_vbr_stackframe;
  wire [3:0] syncreset;
  wire reset;
  wire clkena_lw;
  wire [31:0] tg68_pc;
  wire [31:0] tmp_tg68_pc;
  wire [31:0] tg68_pc_add;
  wire [31:0] pc_dataa;
  wire [31:0] pc_datab;
  wire [31:0] memaddr;
  wire [1:0] state;
  wire [1:0] datatype;
  wire [1:0] set_datatype;
  wire [1:0] exe_datatype;
  wire [1:0] setstate;
  wire setaddrvalue;
  wire addrvalue;
  wire [15:0] opcode;
  wire [15:0] exe_opcode;
  wire [15:0] sndopc;
  wire [31:0] exe_pc  /*verilator public_flat_rd*/ ;
  wire [31:0] last_opc_pc;
  wire [15:0] last_opc_read;
  wire [31:0] reg_qa;
  wire [31:0] reg_qb;
  wire wwrena;
  wire lwrena;
  wire bwrena;
  wire regwrena_now;
  wire [3:0] rf_dest_addr;
  wire [3:0] rf_source_addr;
  wire [3:0] rf_source_addrd;
  wire [31:0] regin;
  wire [3:0] rdindex_a;
  wire [3:0] rdindex_b;
  wire wr_areg;
  wire [31:0] addr;
  wire [31:0] memaddr_reg;
  wire [31:0] memaddr_delta;
  wire [31:0] memaddr_delta_rega;
  wire [31:0] memaddr_delta_regb;
  wire use_base;
  wire [31:0] ea_data;
  wire [31:0] op1out;
  wire [31:0] op2out;
  wire [15:0] op1outbrief;
  wire [31:0] aluout;
  wire [31:0] data_write_tmp;
  wire [31:0] data_write_muxin;
  wire [47:0] data_write_mux;
  wire nextpass;
  wire setnextpass;
  wire setdispbyte;
  wire setdisp;
  wire regdirectsource;
  wire [31:0] addsub_q;
  wire [31:0] briefdata;
  wire [2:0] c_out;
  wire [31:0] memaddr_a;
  wire tg68_pc_brw;
  wire tg68_pc_word;
  wire getbrief;
  wire [15:0] brief;
  wire data_is_source;
  wire store_in_tmp;
  wire write_back;
  wire exec_write_back;
  wire setstackaddr;
  wire writepc;
  wire writepcbig;
  wire set_writepcbig;
  wire writepcnext;
  wire setopcode;
  wire decodeopc  /*verilator public_flat_rd*/ ;
  wire execopc;
  wire execopc_alu;
  wire setexecopc;
  wire endopc;
  wire setendopc;
  wire [7:0] flags /*verilator public_flat_rd*/ ;
  wire [7:0] flagssr /*verilator public_flat_rd*/ ;
  wire [7:0] srin;
  wire exec_direct;
  wire exec_tas;
  wire set_exec_tas;
  wire exe_condition;
  wire ea_only;
  wire source_areg;
  wire source_lowbits;
  wire source_ldrlbits;
  wire source_ldrmbits;
  wire source_2ndhbits;
  wire source_2ndmbits;
  wire source_2ndlbits;
  wire dest_areg;
  wire dest_ldrareg;
  wire dest_ldrhbits;
  wire dest_ldrlbits;
  wire dest_2ndhbits;
  wire dest_2ndlbits;
  wire dest_hbits;
  wire [1:0] rot_bits;
  wire [1:0] set_rot_bits;
  wire [5:0] rot_cnt;
  wire [5:0] set_rot_cnt;
  wire movem_actiond;
  wire [3:0] movem_regaddr;
  wire [3:0] movem_mux;
  wire movem_presub;
  wire movem_run;
  wire set_direct_data;
  wire use_direct_data;
  wire direct_data;
  wire set_v_flag;
  wire set_vectoraddr;
  wire writesr;
  wire trap_berr;
  wire trap_illegal /*verilator public_flat_rd*/ ;
  wire trap_addr_error;
  wire trap_priv;
  wire trap_trace;
  wire trap_1010;
  wire trap_1111;
  wire trap_trap;
  wire trap_trapv;
  wire trap_interrupt;
  wire trapmake;
  wire trapd;
  wire [7:0] trap_sr;
  wire make_trace;
  wire make_berr;
  wire usestackframe2;
  wire set_stop;
  wire stop;
  wire [31:0] trap_vector;
  wire [31:0] trap_vector_vbr;
  wire [31:0] usp;
  wire [2:0] ipl_nr;
  wire [2:0] ripl_nr;
  wire [7:0] ipl_vec;
  wire interrupt;
  wire setinterrupt;
  wire svmode;
  wire presvmode;
  wire suppress_base;
  wire set_suppress_base;
  wire set_z_error;
  wire z_error;
  wire ea_build_now;
  wire build_logical;
  wire build_bcd;
  wire [31:0] data_read;
  wire [7:0] bf_ext_in;
  wire [7:0] bf_ext_out;
  wire long_start;
  wire long_start_alu;
  wire non_aligned;
  wire check_aligned;
  wire long_done;
  wire [5:0] memmask;
  wire [5:0] set_memmask;
  wire [3:0] memread;
  wire [5:0] wbmemmask;
  wire [5:0] memmaskmux;
  wire oddout;
  wire set_oddout;
  wire pcbase;
  wire set_pcbase;
  wire [31:0] last_data_read;
  wire [31:0] last_data_in;
  wire [5:0] bf_offset;
  wire [5:0] bf_width;
  wire [5:0] bf_bhits;
  wire [5:0] bf_shift;
  wire [5:0] alu_width;
  wire [5:0] alu_bf_shift;
  wire [5:0] bf_loffset;
  wire [31:0] bf_full_offset;
  wire [31:0] alu_bf_ffo_offset;
  wire [5:0] alu_bf_loffset;
  wire [31:0] movec_data;
  wire [31:0] vbr;
  wire [3:0] cacr;
  wire [2:0] dfc;
  wire [2:0] sfc;
  wire [88:0] set;
  wire [88:0] set_exec;
  wire [88:0] exec;
  wire [6:0] micro_state;
  wire [6:0] next_micro_state;
  wire [15:0] n34_o;
  wire [15:0] n35_o;
  wire [7:0] alu_n36;
  wire [4:0] n37_o;
  wire alu_n38;
  wire [7:0] alu_n39;
  wire [2:0] alu_n40;
  wire [31:0] alu_n41;
  wire [31:0] alu_n42;
  wire [7:0] alu_bf_ext_out;
  wire alu_set_v_flag;
  wire [7:0] alu_flags;
  wire [2:0] alu_c_out;
  wire [31:0] alu_addsub_q;
  wire [31:0] alu_aluout;
  wire n55_o;
  wire n56_o;
  wire n57_o;
  wire n58_o;
  wire n59_o;
  wire n60_o;
  wire [1:0] n63_o;
  wire n65_o;
  wire [1:0] n66_o;
  wire n68_o;
  wire n69_o;
  wire n72_o;
  wire n77_o;
  wire n78_o;
  wire n81_o;
  wire n82_o;
  wire n84_o;
  wire [5:0] n85_o;
  wire [4:0] n86_o;
  wire [5:0] n88_o;
  wire n89_o;
  wire n90_o;
  wire n92_o;
  wire n93_o;
  wire n94_o;
  wire n97_o;
  wire n98_o;
  wire n102_o;
  wire [2:0] n104_o;
  wire [3:0] n106_o;
  wire n107_o;
  wire n108_o;
  wire n118_o;
  wire n120_o;
  wire n122_o;
  wire n125_o;
  wire n130_o;
  wire n131_o;
  wire [15:0] n132_o;
  wire [31:0] n133_o;
  wire [23:0] n134_o;
  wire [7:0] n135_o;
  wire [31:0] n136_o;
  wire n138_o;
  wire [1:0] n139_o;
  wire n141_o;
  wire n142_o;
  wire n143_o;
  wire n144_o;
  wire n145_o;
  wire n146_o;
  wire n147_o;
  wire n148_o;
  wire n149_o;
  wire n150_o;
  wire n151_o;
  wire n152_o;
  wire n153_o;
  wire n154_o;
  wire n155_o;
  wire n156_o;
  wire n157_o;
  wire n158_o;
  wire n159_o;
  wire n160_o;
  wire [3:0] n161_o;
  wire [3:0] n162_o;
  wire [3:0] n163_o;
  wire [3:0] n164_o;
  wire [15:0] n165_o;
  wire [15:0] n166_o;
  wire [15:0] n167_o;
  wire [15:0] n168_o;
  wire [15:0] n169_o;
  wire [15:0] n170_o;
  wire [15:0] n171_o;
  wire [15:0] n172_o;
  wire n175_o;
  wire n176_o;
  wire n177_o;
  wire n178_o;
  wire [7:0] n179_o;
  wire [7:0] n180_o;
  wire [7:0] n181_o;
  wire n184_o;
  wire n185_o;
  wire n186_o;
  wire n187_o;
  wire n188_o;
  wire n189_o;
  wire n190_o;
  wire n191_o;
  wire n192_o;
  wire n193_o;
  wire n194_o;
  wire n195_o;
  wire n196_o;
  wire n197_o;
  wire n198_o;
  wire n199_o;
  wire n200_o;
  wire n201_o;
  wire n202_o;
  wire n203_o;
  wire n204_o;
  wire n205_o;
  wire n206_o;
  wire n207_o;
  wire n208_o;
  wire n209_o;
  wire n210_o;
  wire n211_o;
  wire [3:0] n212_o;
  wire [3:0] n213_o;
  wire [3:0] n214_o;
  wire [3:0] n215_o;
  wire [15:0] n216_o;
  wire [15:0] n217_o;
  wire [15:0] n218_o;
  wire [15:0] n219_o;
  wire [15:0] n220_o;
  wire [31:0] n221_o;
  wire [31:0] n222_o;
  wire [15:0] n223_o;
  wire [31:0] n224_o;
  wire n225_o;
  wire [31:0] n226_o;
  wire [31:0] n228_o;
  wire [31:0] n229_o;
  wire n233_o;
  wire n234_o;
  wire n235_o;
  wire n236_o;
  wire n240_o;
  wire [31:0] n241_o;
  wire n242_o;
  wire n243_o;
  wire [15:0] n245_o;
  wire [47:0] n246_o;
  wire [39:0] n247_o;
  wire [47:0] n249_o;
  wire [47:0] n250_o;
  wire n251_o;
  wire n252_o;
  wire [15:0] n253_o;
  wire n254_o;
  wire n255_o;
  wire [15:0] n256_o;
  wire [1:0] n257_o;
  wire n259_o;
  wire [7:0] n260_o;
  wire [7:0] n261_o;
  wire [15:0] n262_o;
  wire [1:0] n263_o;
  wire n265_o;
  wire [7:0] n266_o;
  wire [7:0] n267_o;
  wire [15:0] n268_o;
  wire [15:0] n269_o;
  wire [15:0] n270_o;
  wire [15:0] n271_o;
  wire [15:0] n272_o;
  wire [15:0] n273_o;
  wire n274_o;
  wire [7:0] n275_o;
  wire [7:0] n276_o;
  wire [15:0] n277_o;
  wire [15:0] n278_o;
  wire n291_o;
  wire n299_o;
  wire n302_o;
  wire n306_o;
  wire n316_o;
  wire n317_o;
  wire n318_o;
  wire n319_o;
  wire n320_o;
  wire [7:0] n325_o;
  wire [7:0] n326_o;
  wire [7:0] n327_o;
  wire [7:0] n328_o;
  wire [7:0] n329_o;
  wire [7:0] n330_o;
  wire [7:0] n331_o;
  wire [7:0] n332_o;
  wire [7:0] n333_o;
  wire [7:0] n334_o;
  wire [7:0] n335_o;
  wire [15:0] n336_o;
  wire [15:0] n337_o;
  wire [15:0] n338_o;
  wire [15:0] n339_o;
  wire [15:0] n340_o;
  wire [15:0] n341_o;
  wire [15:0] n342_o;
  wire [15:0] n343_o;
  wire [15:0] n344_o;
  wire [7:0] n345_o;
  wire [7:0] n346_o;
  wire [7:0] n347_o;
  wire [7:0] n348_o;
  wire [7:0] n349_o;
  wire [7:0] n350_o;
  wire [7:0] n351_o;
  wire [7:0] n352_o;
  wire [7:0] n353_o;
  wire n354_o;
  wire [15:0] n355_o;
  wire [15:0] n356_o;
  wire n357_o;
  wire n358_o;
  wire n359_o;
  wire n360_o;
  wire n361_o;
  wire n362_o;
  wire n364_o;
  wire n365_o;
  wire n368_o;
  wire n370_o;
  wire [1:0] n371_o;
  reg n374_o;
  reg n377_o;
  wire n380_o;
  wire n382_o;
  wire n384_o;
  wire n386_o;
  wire n388_o;
  wire n390_o;
  wire n392_o;
  wire n395_o;
  wire n398_o;
  wire n403_o;
  wire n404_o;
  wire [3:0] n405_o;
  wire n406_o;
  wire [2:0] n407_o;
  wire [3:0] n409_o;
  wire [2:0] n410_o;
  wire [3:0] n411_o;
  wire [3:0] n412_o;
  wire [2:0] n413_o;
  wire [3:0] n415_o;
  wire [2:0] n416_o;
  wire [3:0] n418_o;
  wire [2:0] n419_o;
  wire [3:0] n420_o;
  wire [2:0] n421_o;
  wire n423_o;
  wire n424_o;
  wire [2:0] n425_o;
  wire [3:0] n426_o;
  wire [2:0] n427_o;
  wire [3:0] n429_o;
  wire [3:0] n430_o;
  wire [3:0] n431_o;
  wire [3:0] n433_o;
  wire [3:0] n434_o;
  wire [3:0] n435_o;
  wire [3:0] n436_o;
  wire [3:0] n437_o;
  wire [3:0] n438_o;
  wire [3:0] n439_o;
  wire [3:0] n440_o;
  wire n444_o;
  wire n445_o;
  wire n446_o;
  wire [3:0] n448_o;
  wire [3:0] n449_o;
  wire [2:0] n450_o;
  wire [3:0] n452_o;
  wire [2:0] n453_o;
  wire [3:0] n455_o;
  wire [2:0] n456_o;
  wire [3:0] n458_o;
  wire [2:0] n459_o;
  wire [3:0] n461_o;
  wire [2:0] n462_o;
  wire [3:0] n464_o;
  wire [2:0] n465_o;
  wire [3:0] n466_o;
  wire n467_o;
  wire [2:0] n468_o;
  wire [3:0] n469_o;
  wire [3:0] n471_o;
  wire [3:0] n472_o;
  wire [3:0] n473_o;
  wire [3:0] n474_o;
  wire [3:0] n475_o;
  wire [3:0] n476_o;
  wire [3:0] n477_o;
  wire [3:0] n478_o;
  wire n482_o;
  wire n483_o;
  wire n484_o;
  wire n485_o;
  wire n486_o;
  wire n487_o;
  wire n488_o;
  wire n489_o;
  wire n490_o;
  wire [31:0] n491_o;
  wire [31:0] n492_o;
  wire [31:0] n494_o;
  wire [15:0] n498_o;
  wire n499_o;
  wire n500_o;
  wire n501_o;
  wire n502_o;
  wire n503_o;
  wire n504_o;
  wire n505_o;
  wire n506_o;
  wire n507_o;
  wire n508_o;
  wire n509_o;
  wire n510_o;
  wire n511_o;
  wire n512_o;
  wire n513_o;
  wire n514_o;
  wire [3:0] n515_o;
  wire [3:0] n516_o;
  wire [3:0] n517_o;
  wire [3:0] n518_o;
  wire [15:0] n519_o;
  wire n520_o;
  localparam [15:0] n521_o = 16'b1111111111111111;
  wire n522_o;
  wire n523_o;
  wire n524_o;
  wire n525_o;
  wire n526_o;
  wire n527_o;
  wire n528_o;
  wire n529_o;
  wire n530_o;
  wire n531_o;
  wire n532_o;
  wire [7:0] n533_o;
  wire n534_o;
  wire n535_o;
  wire n536_o;
  wire n537_o;
  wire n538_o;
  wire n539_o;
  wire n540_o;
  wire n541_o;
  wire [3:0] n542_o;
  wire [3:0] n543_o;
  wire [7:0] n544_o;
  wire n545_o;
  wire [2:0] n546_o;
  wire [2:0] n547_o;
  wire n549_o;
  wire n552_o;
  wire n555_o;
  wire n556_o;
  wire n557_o;
  wire n558_o;
  wire [15:0] n559_o;
  wire [15:0] n560_o;
  wire [15:0] n561_o;
  wire [15:0] n562_o;
  wire [15:0] n563_o;
  wire [31:0] n564_o;
  wire [15:0] n565_o;
  wire [15:0] n566_o;
  wire [15:0] n567_o;
  wire [15:0] n568_o;
  wire [15:0] n569_o;
  wire [31:0] n570_o;
  wire [31:0] n571_o;
  wire [31:0] n572_o;
  wire [15:0] n575_o;
  wire [15:0] n576_o;
  wire n577_o;
  wire n578_o;
  wire n579_o;
  wire n580_o;
  wire n581_o;
  wire n582_o;
  wire n583_o;
  wire n584_o;
  wire n585_o;
  wire n586_o;
  wire n587_o;
  wire n588_o;
  wire n589_o;
  wire n590_o;
  wire n591_o;
  wire n592_o;
  wire n593_o;
  wire n594_o;
  wire n595_o;
  wire n596_o;
  wire n597_o;
  wire n598_o;
  wire n599_o;
  wire n600_o;
  wire n601_o;
  wire [3:0] n602_o;
  wire [3:0] n603_o;
  wire [3:0] n604_o;
  wire [3:0] n605_o;
  wire [3:0] n606_o;
  wire [3:0] n607_o;
  wire [15:0] n608_o;
  wire [7:0] n609_o;
  wire [23:0] n610_o;
  wire [7:0] n611_o;
  wire [7:0] n612_o;
  wire [7:0] n613_o;
  wire [7:0] n614_o;
  wire [7:0] n615_o;
  wire [7:0] n616_o;
  wire [7:0] n617_o;
  wire [23:0] n618_o;
  wire [23:0] n619_o;
  wire [7:0] n620_o;
  wire [7:0] n621_o;
  wire [7:0] n622_o;
  wire [7:0] n623_o;
  wire [7:0] n624_o;
  wire [7:0] n625_o;
  wire [7:0] n626_o;
  wire n631_o;
  wire n633_o;
  wire n634_o;
  wire n635_o;
  wire n637_o;
  wire n639_o;
  wire n642_o;
  wire n644_o;
  wire n646_o;
  wire n647_o;
  wire n649_o;
  wire n650_o;
  wire n652_o;
  wire n654_o;
  wire n655_o;
  wire n656_o;
  wire n658_o;
  wire n660_o;
  wire n661_o;
  wire n663_o;
  wire n665_o;
  wire n667_o;
  wire n668_o;
  wire n670_o;
  wire n672_o;
  wire n673_o;
  wire n674_o;
  wire n675_o;
  wire n676_o;
  wire n677_o;
  wire n679_o;
  wire n680_o;
  wire n681_o;
  wire [31:0] n682_o;
  wire [31:0] n683_o;
  wire [31:0] n684_o;
  wire n685_o;
  wire n687_o;
  wire n689_o;
  wire n690_o;
  wire n692_o;
  wire n693_o;
  wire n694_o;
  wire n695_o;
  wire n696_o;
  wire n698_o;
  wire [11:0] n699_o;
  wire [15:0] n701_o;
  wire n702_o;
  wire [11:0] n703_o;
  wire [15:0] n705_o;
  wire n706_o;
  wire n707_o;
  wire n708_o;
  wire n709_o;
  wire [11:0] n710_o;
  wire [15:0] n712_o;
  wire n713_o;
  wire n714_o;
  wire n715_o;
  wire n716_o;
  wire [15:0] n717_o;
  wire n718_o;
  wire [15:0] n719_o;
  wire n720_o;
  wire n721_o;
  wire n722_o;
  wire n723_o;
  wire n724_o;
  wire n726_o;
  wire n727_o;
  wire n728_o;
  wire [23:0] n729_o;
  wire [23:0] n730_o;
  wire [23:0] n731_o;
  wire [7:0] n732_o;
  wire n733_o;
  wire [15:0] n734_o;
  wire [15:0] n735_o;
  wire [15:0] n736_o;
  wire [15:0] n737_o;
  wire [15:0] n738_o;
  wire [15:0] n739_o;
  wire [15:0] n740_o;
  wire [31:0] n741_o;
  wire [31:0] n742_o;
  wire [15:0] n743_o;
  wire [15:0] n744_o;
  wire [15:0] n745_o;
  wire [15:0] n746_o;
  wire [15:0] n747_o;
  wire [31:0] n748_o;
  wire [31:0] n749_o;
  wire [31:0] n750_o;
  wire [31:0] n751_o;
  wire [31:0] n752_o;
  wire [31:0] n753_o;
  wire [31:0] n754_o;
  wire [15:0] n755_o;
  wire [15:0] n756_o;
  wire [15:0] n757_o;
  wire [15:0] n758_o;
  wire [15:0] n759_o;
  wire n760_o;
  wire [31:0] n761_o;
  wire [31:0] n762_o;
  wire n763_o;
  wire n766_o;
  wire [31:0] n768_o;
  wire n769_o;
  wire n771_o;
  wire [31:0] n772_o;
  wire n773_o;
  wire n775_o;
  wire [31:0] n776_o;
  wire n777_o;
  wire n779_o;
  wire [31:0] n781_o;
  wire [31:0] n782_o;
  wire n783_o;
  wire n784_o;
  wire n785_o;
  wire n786_o;
  wire n787_o;
  wire n788_o;
  wire n789_o;
  wire [31:0] n790_o;
  wire [31:0] n791_o;
  wire n793_o;
  wire n795_o;
  wire n796_o;
  wire n798_o;
  wire n800_o;
  wire n801_o;
  wire n803_o;
  wire n816_o;
  wire [15:0] n817_o;
  wire n818_o;
  wire n819_o;
  wire n820_o;
  wire n821_o;
  wire n822_o;
  wire n823_o;
  wire n824_o;
  wire n825_o;
  wire n826_o;
  wire n827_o;
  wire n828_o;
  wire n829_o;
  wire n830_o;
  wire n831_o;
  wire n832_o;
  wire n833_o;
  wire [3:0] n834_o;
  wire [3:0] n835_o;
  wire [3:0] n836_o;
  wire [3:0] n837_o;
  wire [15:0] n838_o;
  wire [15:0] n839_o;
  wire [15:0] n840_o;
  wire [31:0] n841_o;
  wire n842_o;
  wire n844_o;
  wire n846_o;
  wire [1:0] n847_o;
  wire [15:0] n848_o;
  wire [31:0] n849_o;
  wire n851_o;
  wire [14:0] n852_o;
  wire [15:0] n853_o;
  wire [30:0] n854_o;
  wire [31:0] n856_o;
  wire n858_o;
  wire [13:0] n859_o;
  wire [15:0] n860_o;
  wire [29:0] n861_o;
  wire [31:0] n863_o;
  wire n865_o;
  wire [12:0] n866_o;
  wire [15:0] n867_o;
  wire [28:0] n868_o;
  wire [31:0] n870_o;
  wire n872_o;
  wire [3:0] n873_o;
  reg [31:0] n874_o;
  wire [31:0] n875_o;
  wire [9:0] n882_o;
  wire [9:0] n883_o;
  wire [9:0] n885_o;
  wire [9:0] n887_o;
  wire [9:0] n889_o;
  wire n890_o;
  wire [9:0] n892_o;
  wire [9:0] n894_o;
  wire [9:0] n896_o;
  wire [9:0] n898_o;
  wire [9:0] n900_o;
  wire [9:0] n902_o;
  wire [3:0] n903_o;
  wire [7:0] n905_o;
  wire [9:0] n907_o;
  wire [9:0] n908_o;
  wire n909_o;
  wire [9:0] n911_o;
  wire [9:0] n912_o;
  wire [31:0] n913_o;
  wire [31:0] n916_o;
  wire [31:0] n917_o;
  wire n919_o;
  wire n920_o;
  wire n921_o;
  wire [2:0] n922_o;
  wire n923_o;
  wire n924_o;
  wire n925_o;
  wire n926_o;
  wire n927_o;
  wire n928_o;
  wire n929_o;
  wire n930_o;
  wire [3:0] n931_o;
  wire [3:0] n932_o;
  wire [7:0] n933_o;
  wire n934_o;
  wire n935_o;
  wire n936_o;
  wire n937_o;
  wire n938_o;
  wire n939_o;
  wire n940_o;
  wire n941_o;
  wire n942_o;
  wire n943_o;
  wire n944_o;
  wire n945_o;
  wire n946_o;
  wire n947_o;
  wire n948_o;
  wire n949_o;
  wire [3:0] n950_o;
  wire [3:0] n951_o;
  wire [3:0] n952_o;
  wire [3:0] n953_o;
  wire [15:0] n954_o;
  wire n955_o;
  wire [31:0] n956_o;
  wire [7:0] n957_o;
  wire [7:0] n958_o;
  wire [7:0] n959_o;
  wire [23:0] n960_o;
  wire [23:0] n961_o;
  wire [23:0] n962_o;
  wire [31:0] n963_o;
  wire [31:0] n964_o;
  wire n965_o;
  wire n966_o;
  wire n969_o;
  wire n970_o;
  wire n971_o;
  wire n972_o;
  wire [4:0] n975_o;
  wire [4:0] n976_o;
  wire [3:0] n978_o;
  wire [4:0] n980_o;
  wire [4:0] n981_o;
  wire [4:0] n982_o;
  wire [4:0] n983_o;
  wire [4:0] n984_o;
  wire [26:0] n985_o;
  wire [26:0] n986_o;
  wire [26:0] n987_o;
  wire n989_o;
  wire n991_o;
  wire n992_o;
  wire n993_o;
  wire n994_o;
  wire n996_o;
  wire n997_o;
  wire n998_o;
  wire n999_o;
  wire n1000_o;
  wire n1001_o;
  wire n1002_o;
  wire n1004_o;
  wire n1005_o;
  wire n1006_o;
  wire n1008_o;
  wire n1009_o;
  wire n1010_o;
  wire n1011_o;
  wire n1012_o;
  wire n1015_o;
  wire [31:0] n1016_o;
  wire n1018_o;
  wire [31:0] n1019_o;
  wire [31:0] n1021_o;
  wire n1023_o;
  wire [31:0] n1024_o;
  wire [31:0] n1026_o;
  wire n1028_o;
  wire [31:0] n1029_o;
  wire [31:0] n1031_o;
  wire n1033_o;
  wire [31:0] n1034_o;
  wire [31:0] n1036_o;
  wire n1038_o;
  wire [31:0] n1039_o;
  wire [31:0] n1041_o;
  wire n1043_o;
  wire [31:0] n1044_o;
  wire [31:0] n1046_o;
  wire n1048_o;
  wire [31:0] n1049_o;
  wire [31:0] n1051_o;
  wire n1054_o;
  wire n1056_o;
  wire n1057_o;
  wire n1058_o;
  wire n1059_o;
  wire n1060_o;
  wire n1062_o;
  wire n1063_o;
  wire [31:0] n1072_o;
  wire [31:0] n1073_o;
  wire [31:0] n1074_o;
  wire n1075_o;
  wire [31:0] n1077_o;
  wire [31:0] n1081_o;
  localparam [2:0] n1082_o = 3'b000;
  wire n1083_o;
  wire n1084_o;
  wire n1085_o;
  wire n1086_o;
  wire n1087_o;
  wire [3:0] n1088_o;
  wire n1089_o;
  wire n1090_o;
  wire n1091_o;
  wire n1092_o;
  wire n1093_o;
  wire n1094_o;
  wire n1095_o;
  wire n1096_o;
  wire [3:0] n1097_o;
  wire [3:0] n1098_o;
  wire [7:0] n1099_o;
  wire n1100_o;
  wire n1101_o;
  wire n1102_o;
  wire n1103_o;
  wire n1104_o;
  wire n1105_o;
  wire n1106_o;
  wire n1107_o;
  wire n1108_o;
  wire n1109_o;
  wire n1110_o;
  wire n1111_o;
  wire n1112_o;
  wire n1113_o;
  wire n1114_o;
  wire n1115_o;
  wire [3:0] n1116_o;
  wire [3:0] n1117_o;
  wire [3:0] n1118_o;
  wire [3:0] n1119_o;
  wire [15:0] n1120_o;
  localparam [1:0] n1121_o = 2'b11;
  wire n1124_o;
  wire n1125_o;
  wire n1129_o;
  wire n1130_o;
  wire n1131_o;
  wire n1132_o;
  wire n1133_o;
  wire n1134_o;
  wire n1135_o;
  wire n1136_o;
  wire n1137_o;
  wire n1138_o;
  wire n1139_o;
  wire n1140_o;
  wire n1141_o;
  wire n1142_o;
  wire n1143_o;
  wire n1144_o;
  wire n1146_o;
  wire n1148_o;
  wire n1150_o;
  wire n1151_o;
  wire n1152_o;
  wire n1153_o;
  wire [2:0] n1154_o;
  wire n1155_o;
  wire n1156_o;
  wire [1:0] n1157_o;
  wire n1158_o;
  wire n1159_o;
  wire n1160_o;
  wire [1:0] n1161_o;
  wire [1:0] n1162_o;
  wire [7:0] n1166_o;
  wire [7:0] n1167_o;
  wire [7:0] n1168_o;
  wire [23:0] n1169_o;
  wire [23:0] n1170_o;
  wire [23:0] n1171_o;
  wire [31:0] n1172_o;
  wire [31:0] n1173_o;
  wire [31:0] n1174_o;
  wire [31:0] n1175_o;
  wire n1177_o;
  wire n1179_o;
  wire n1180_o;
  wire n1181_o;
  wire n1182_o;
  wire n1183_o;
  wire n1185_o;
  wire n1186_o;
  wire n1187_o;
  wire n1189_o;
  wire n1190_o;
  wire n1191_o;
  wire n1192_o;
  wire n1193_o;
  wire [2:0] n1194_o;
  wire n1195_o;
  wire n1197_o;
  wire n1198_o;
  wire n1199_o;
  wire n1200_o;
  wire n1201_o;
  wire n1204_o;
  wire n1206_o;
  wire n1209_o;
  wire n1211_o;
  wire n1215_o;
  wire n1218_o;
  wire n1221_o;
  wire n1223_o;
  wire n1224_o;
  wire n1225_o;
  wire n1226_o;
  wire n1227_o;
  wire n1229_o;
  wire n1230_o;
  wire n1231_o;
  wire n1232_o;
  wire n1233_o;
  wire n1236_o;
  wire [2:0] n1238_o;
  wire [3:0] n1240_o;
  wire [5:0] n1242_o;
  wire [1:0] n1243_o;
  wire [1:0] n1244_o;
  wire [3:0] n1245_o;
  wire n1246_o;
  wire n1247_o;
  wire n1249_o;
  wire n1250_o;
  wire n1251_o;
  wire n1252_o;
  wire [31:0] n1253_o;
  wire [31:0] n1254_o;
  wire [31:0] n1255_o;
  wire [31:0] n1256_o;
  wire [5:0] n1257_o;
  wire [3:0] n1258_o;
  wire n1259_o;
  wire n1260_o;
  wire n1262_o;
  wire n1263_o;
  wire n1264_o;
  wire n1265_o;
  wire [7:0] n1267_o;
  wire n1270_o;
  wire n1273_o;
  wire [2:0] n1274_o;
  wire [7:0] n1275_o;
  wire n1277_o;
  wire n1281_o;
  wire n1284_o;
  wire [2:0] n1286_o;
  wire [7:0] n1287_o;
  wire n1288_o;
  wire n1289_o;
  wire n1290_o;
  wire n1292_o;
  wire [2:0] n1293_o;
  wire [7:0] n1294_o;
  wire n1296_o;
  wire n1297_o;
  wire n1298_o;
  wire [7:0] n1299_o;
  wire [7:0] n1300_o;
  wire n1302_o;
  wire [15:0] n1303_o;
  wire [31:0] n1304_o;
  wire [15:0] n1305_o;
  wire [7:0] n1306_o;
  wire n1308_o;
  wire [7:0] n1309_o;
  wire n1311_o;
  wire n1312_o;
  wire n1313_o;
  wire n1315_o;
  wire n1317_o;
  wire n1319_o;
  wire n1321_o;
  wire n1323_o;
  wire n1324_o;
  wire [31:0] n1325_o;
  wire [31:0] n1326_o;
  wire [31:0] n1328_o;
  wire [5:0] n1329_o;
  wire [5:0] n1330_o;
  wire [31:0] n1331_o;
  wire [5:0] n1332_o;
  wire n1333_o;
  wire n1334_o;
  wire n1335_o;
  wire n1336_o;
  wire n1337_o;
  wire n1338_o;
  wire n1339_o;
  wire n1340_o;
  wire n1341_o;
  wire n1342_o;
  wire n1343_o;
  wire [1:0] n1345_o;
  wire [1:0] n1346_o;
  wire n1348_o;
  wire n1350_o;
  wire n1351_o;
  wire n1352_o;
  wire n1353_o;
  wire n1355_o;
  wire n1357_o;
  wire n1359_o;
  wire n1360_o;
  wire n1361_o;
  wire n1362_o;
  wire n1364_o;
  wire n1365_o;
  wire n1367_o;
  wire n1368_o;
  wire n1369_o;
  wire n1370_o;
  wire n1371_o;
  wire n1372_o;
  wire n1373_o;
  wire n1374_o;
  wire n1377_o;
  wire n1378_o;
  wire n1379_o;
  wire n1381_o;
  wire n1382_o;
  wire n1383_o;
  wire n1384_o;
  wire n1387_o;
  wire [5:0] n1390_o;
  wire [5:0] n1393_o;
  wire n1395_o;
  wire [5:0] n1397_o;
  wire [5:0] n1399_o;
  wire n1401_o;
  wire [5:0] n1402_o;
  wire [5:0] n1403_o;
  wire n1404_o;
  wire [5:0] n1406_o;
  wire [5:0] n1408_o;
  wire n1409_o;
  wire [1:0] n1410_o;
  wire [1:0] n1412_o;
  wire n1414_o;
  wire [5:0] n1415_o;
  wire [5:0] n1416_o;
  wire n1417_o;
  wire [1:0] n1418_o;
  wire [1:0] n1420_o;
  wire n1422_o;
  wire [5:0] n1424_o;
  wire [5:0] n1425_o;
  wire n1426_o;
  wire n1427_o;
  wire n1429_o;
  wire [1:0] n1430_o;
  wire n1431_o;
  wire n1432_o;
  wire n1434_o;
  wire n1435_o;
  wire [5:0] n1436_o;
  wire n1437_o;
  wire n1438_o;
  wire n1439_o;
  wire n1440_o;
  wire n1442_o;
  wire n1444_o;
  wire n1445_o;
  wire [15:0] n1446_o;
  wire [15:0] n1447_o;
  wire [15:0] n1448_o;
  wire n1449_o;
  wire n1450_o;
  wire n1452_o;
  wire [15:0] n1453_o;
  wire [15:0] n1454_o;
  wire [31:0] n1455_o;
  wire n1456_o;
  wire n1457_o;
  wire n1459_o;
  wire [15:0] n1461_o;
  wire n1463_o;
  wire [15:0] n1464_o;
  wire [31:0] n1465_o;
  wire n1467_o;
  wire n1468_o;
  wire [7:0] n1469_o;
  wire [1:0] n1470_o;
  wire [1:0] n1471_o;
  wire [1:0] n1472_o;
  wire [1:0] n1473_o;
  wire n1474_o;
  wire [15:0] n1475_o;
  wire [15:0] n1476_o;
  wire n1477_o;
  wire n1478_o;
  wire n1479_o;
  wire n1480_o;
  wire n1481_o;
  wire n1482_o;
  wire n1483_o;
  wire n1484_o;
  wire n1485_o;
  wire n1486_o;
  wire n1487_o;
  wire n1488_o;
  wire n1489_o;
  wire n1490_o;
  wire n1491_o;
  wire n1492_o;
  wire n1493_o;
  wire n1494_o;
  wire n1495_o;
  wire n1496_o;
  wire [7:0] n1497_o;
  wire n1498_o;
  wire n1499_o;
  wire [5:0] n1500_o;
  wire [3:0] n1502_o;
  wire [5:0] n1503_o;
  wire n1504_o;
  wire n1505_o;
  wire n1506_o;
  wire n1507_o;
  wire n1508_o;
  wire [1:0] n1509_o;
  wire [1:0] n1510_o;
  wire [31:0] n1512_o;
  wire [1:0] n1514_o;
  wire [1:0] n1515_o;
  wire n1517_o;
  wire [15:0] n1519_o;
  wire [15:0] n1520_o;
  wire [31:0] n1521_o;
  wire [31:0] n1522_o;
  wire [15:0] n1524_o;
  wire n1525_o;
  wire n1527_o;
  wire [15:0] n1528_o;
  wire n1530_o;
  wire n1532_o;
  wire n1534_o;
  wire n1536_o;
  wire n1538_o;
  wire [1:0] n1539_o;
  wire [5:0] n1541_o;
  wire n1543_o;
  wire n1545_o;
  wire n1547_o;
  wire [7:0] n1548_o;
  wire n1550_o;
  wire n1552_o;
  wire [2:0] n1553_o;
  wire [7:0] n1554_o;
  wire n1556_o;
  wire n1558_o;
  wire [5:0] n1560_o;
  wire [3:0] n1561_o;
  wire [5:0] n1562_o;
  wire n1563_o;
  wire [5:0] n1564_o;
  wire [5:0] n1565_o;
  wire [31:0] n1566_o;
  wire [5:0] n1567_o;
  wire n1608_o;
  wire n1609_o;
  wire n1610_o;
  wire n1611_o;
  wire n1612_o;
  wire n1614_o;
  wire n1615_o;
  wire n1617_o;
  wire n1618_o;
  wire n1619_o;
  wire n1620_o;
  wire n1623_o;
  wire n1624_o;
  wire n1625_o;
  wire [1:0] n1626_o;
  wire n1627_o;
  wire n1628_o;
  wire n1629_o;
  wire [35:0] n1630_o;
  wire [47:0] n1631_o;
  wire [88:0] n1632_o;
  wire n1633_o;
  wire n1634_o;
  wire n1635_o;
  wire n1636_o;
  wire n1637_o;
  wire [84:0] n1639_o;
  wire n1640_o;
  wire n1641_o;
  wire n1642_o;
  wire n1643_o;
  wire n1644_o;
  wire [1:0] n1645_o;
  wire n1647_o;
  wire [88:0] n1649_o;
  wire [88:0] n1650_o;
  wire n1652_o;
  wire n1653_o;
  wire [16:0] n1654_o;
  wire [16:0] n1655_o;
  wire [16:0] n1656_o;
  wire [70:0] n1657_o;
  wire [70:0] n1658_o;
  wire [70:0] n1659_o;
  wire [88:0] n1661_o;
  wire n1669_o;
  wire [4:0] n1670_o;
  wire [5:0] n1672_o;
  wire [4:0] n1673_o;
  wire [5:0] n1675_o;
  wire n1677_o;
  wire [4:0] n1678_o;
  localparam [31:0] n1679_o = 32'b00000000000000000000000000000000;
  wire [26:0] n1680_o;
  wire [31:0] n1681_o;
  wire [31:0] n1682_o;
  wire n1684_o;
  wire [4:0] n1685_o;
  wire [4:0] n1687_o;
  wire [4:0] n1688_o;
  wire [4:0] n1690_o;
  wire [4:0] n1691_o;
  wire [5:0] n1692_o;
  wire n1693_o;
  wire n1694_o;
  wire [2:0] n1695_o;
  wire n1697_o;
  wire [5:0] n1699_o;
  wire [4:0] n1702_o;
  wire [4:0] n1703_o;
  wire [4:0] n1704_o;
  wire [1:0] n1705_o;
  wire n1707_o;
  wire [2:0] n1708_o;
  wire n1710_o;
  wire [5:0] n1712_o;
  wire [5:0] n1714_o;
  wire [4:0] n1717_o;
  wire [4:0] n1718_o;
  wire [4:0] n1719_o;
  wire [2:0] n1720_o;
  wire n1722_o;
  wire [2:0] n1723_o;
  wire [5:0] n1725_o;
  wire [5:0] n1727_o;
  wire [4:0] n1729_o;
  wire [2:0] n1730_o;
  wire [2:0] n1732_o;
  wire [5:0] n1734_o;
  wire [5:0] n1735_o;
  wire [5:0] n1736_o;
  wire [1:0] n1738_o;
  wire [1:0] n1739_o;
  wire [1:0] n1740_o;
  wire [1:0] n1741_o;
  wire n1742_o;
  wire n1743_o;
  wire n1744_o;
  wire [2:0] n1745_o;
  wire [2:0] n1746_o;
  wire [2:0] n1747_o;
  wire [5:0] n1748_o;
  wire [5:0] n1749_o;
  wire [2:0] n1750_o;
  wire n1752_o;
  wire n1754_o;
  wire n1756_o;
  wire n1758_o;
  wire [3:0] n1759_o;
  reg [5:0] n1765_o;
  wire n1767_o;
  wire [5:0] n1769_o;
  wire n1773_o;
  wire [7:0] n1774_o;
  wire [7:0] n1775_o;
  wire n1776_o;
  wire [7:0] n1777_o;
  wire [7:0] n1778_o;
  wire n1779_o;
  wire [7:0] n1780_o;
  wire [7:0] n1781_o;
  wire [7:0] n1782_o;
  wire [7:0] n1783_o;
  wire [7:0] n1784_o;
  wire [7:0] n1785_o;
  wire n1788_o;
  wire n1789_o;
  wire n1790_o;
  wire n1791_o;
  wire n1792_o;
  wire n1793_o;
  wire n1794_o;
  wire n1795_o;
  wire n1796_o;
  wire n1797_o;
  wire n1798_o;
  wire n1800_o;
  wire n1801_o;
  wire n1803_o;
  wire n1804_o;
  wire n1805_o;
  wire n1806_o;
  wire n1807_o;
  wire n1808_o;
  wire n1809_o;
  wire n1810_o;
  wire n1811_o;
  wire n1812_o;
  wire n1814_o;
  wire n1816_o;
  wire n1818_o;
  wire n1819_o;
  wire n1821_o;
  wire n1822_o;
  wire n1823_o;
  wire [4:0] n1825_o;
  wire n1826_o;
  wire [7:0] n1827_o;
  wire n1829_o;
  wire [2:0] n1830_o;
  wire [2:0] n1831_o;
  wire [2:0] n1832_o;
  wire [2:0] n1833_o;
  wire [4:0] n1834_o;
  wire [4:0] n1835_o;
  wire [4:0] n1836_o;
  wire n1837_o;
  wire n1838_o;
  wire n1839_o;
  wire n1840_o;
  wire n1841_o;
  wire n1842_o;
  wire [7:0] n1843_o;
  wire n1846_o;
  wire n1847_o;
  wire n1848_o;
  wire n1851_o;
  wire n1852_o;
  wire n1853_o;
  wire n1854_o;
  wire n1855_o;
  wire n1856_o;
  wire n1857_o;
  wire n1858_o;
  wire n1865_o;
  wire n1866_o;
  wire n1867_o;
  wire n1868_o;
  wire n1869_o;
  wire n1870_o;
  wire [2:0] n1872_o;
  wire [2:0] n1873_o;
  wire [2:0] n1874_o;
  wire n1875_o;
  wire n1876_o;
  wire [7:0] n1877_o;
  wire [7:0] n1878_o;
  wire n1879_o;
  wire n1880_o;
  wire n1881_o;
  wire n1882_o;
  wire [7:0] n1884_o;
  wire n1886_o;
  wire n1888_o;
  wire n1890_o;
  wire [1:0] n1900_o;
  wire n1902_o;
  wire [5:0] n1904_o;
  localparam [5:0] n1905_o = 6'b000001;
  wire [5:0] n1906_o;
  localparam [88:0] n1909_o = 89'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  wire [1:0] n1912_o;
  wire n1914_o;
  wire n1916_o;
  wire [1:0] n1917_o;
  reg [1:0] n1921_o;
  wire n1922_o;
  wire n1924_o;
  wire n1925_o;
  wire n1928_o;
  wire n1929_o;
  wire n1931_o;
  wire n1932_o;
  wire [1:0] n1935_o;
  wire n1938_o;
  wire [1:0] n1940_o;
  wire [6:0] n1943_o;
  wire n1945_o;
  wire n1946_o;
  wire n1947_o;
  wire n1948_o;
  wire n1949_o;
  wire n1950_o;
  wire n1951_o;
  wire [6:0] n1954_o;
  wire [6:0] n1956_o;
  wire n1957_o;
  wire n1959_o;
  wire n1960_o;
  wire n1961_o;
  wire n1963_o;
  wire [1:0] n1965_o;
  wire n1967_o;
  wire n1968_o;
  wire [6:0] n1971_o;
  wire n1973_o;
  wire n1974_o;
  wire n1975_o;
  wire n1976_o;
  wire n1977_o;
  wire [6:0] n1980_o;
  wire n1981_o;
  wire n1983_o;
  wire [1:0] n1985_o;
  wire n1986_o;
  wire [6:0] n1987_o;
  wire n1989_o;
  wire n1990_o;
  wire n1991_o;
  wire n1992_o;
  wire n1994_o;
  wire [1:0] n1996_o;
  wire n1997_o;
  wire n1998_o;
  wire n1999_o;
  wire n2000_o;
  wire n2002_o;
  wire n2003_o;
  wire [1:0] n2006_o;
  wire n2007_o;
  wire [6:0] n2009_o;
  wire n2010_o;
  wire n2015_o;
  wire [1:0] n2017_o;
  wire [1:0] n2018_o;
  wire [1:0] n2019_o;
  wire n2022_o;
  wire n2023_o;
  wire n2024_o;
  wire [1:0] n2026_o;
  wire n2027_o;
  wire n2028_o;
  wire n2029_o;
  wire n2031_o;
  wire n2032_o;
  wire n2035_o;
  wire n2036_o;
  wire n2037_o;
  wire [2:0] n2038_o;
  wire n2040_o;
  wire [2:0] n2042_o;
  wire n2044_o;
  wire n2046_o;
  wire n2047_o;
  wire n2048_o;
  wire n2049_o;
  wire n2051_o;
  wire n2052_o;
  wire [2:0] n2054_o;
  wire n2056_o;
  wire n2058_o;
  wire n2059_o;
  wire n2060_o;
  wire n2061_o;
  wire n2063_o;
  wire n2065_o;
  wire n2066_o;
  wire n2068_o;
  wire n2069_o;
  wire n2071_o;
  wire n2073_o;
  wire [2:0] n2074_o;
  wire n2076_o;
  wire n2079_o;
  wire n2082_o;
  wire n2085_o;
  wire n2087_o;
  wire n2089_o;
  wire n2091_o;
  wire [4:0] n2092_o;
  reg n2095_o;
  reg n2098_o;
  reg n2101_o;
  reg n2105_o;
  reg n2109_o;
  wire n2110_o;
  reg n2111_o;
  reg n2112_o;
  reg [6:0] n2117_o;
  wire n2119_o;
  wire [3:0] n2120_o;
  reg n2123_o;
  reg n2126_o;
  reg n2128_o;
  reg n2130_o;
  reg n2132_o;
  wire n2133_o;
  reg n2134_o;
  wire n2135_o;
  reg n2136_o;
  wire n2137_o;
  reg n2138_o;
  wire n2139_o;
  reg n2140_o;
  wire n2141_o;
  reg n2142_o;
  reg n2143_o;
  reg [6:0] n2146_o;
  wire n2148_o;
  wire n2151_o;
  wire n2154_o;
  wire n2157_o;
  wire n2160_o;
  wire [1:0] n2162_o;
  wire n2163_o;
  wire n2164_o;
  wire [1:0] n2165_o;
  wire [1:0] n2166_o;
  wire n2167_o;
  wire n2168_o;
  wire n2169_o;
  wire n2170_o;
  wire n2171_o;
  wire [1:0] n2177_o;
  wire [1:0] n2178_o;
  wire [10:0] n2179_o;
  wire [6:0] n2180_o;
  wire n2181_o;
  wire n2183_o;
  wire n2184_o;
  wire [3:0] n2185_o;
  wire n2186_o;
  wire [2:0] n2187_o;
  wire n2189_o;
  wire n2190_o;
  wire n2193_o;
  wire n2194_o;
  wire n2198_o;
  wire n2199_o;
  wire n2201_o;
  wire n2203_o;
  wire n2204_o;
  wire n2206_o;
  wire n2207_o;
  wire n2208_o;
  wire n2210_o;
  wire n2211_o;
  wire n2212_o;
  wire [6:0] n2214_o;
  wire n2217_o;
  wire n2218_o;
  wire [2:0] n2219_o;
  wire n2221_o;
  wire n2222_o;
  wire [2:0] n2223_o;
  wire n2225_o;
  wire [5:0] n2226_o;
  wire n2228_o;
  wire n2229_o;
  wire n2230_o;
  wire n2231_o;
  wire n2232_o;
  wire [6:0] n2233_o;
  wire n2235_o;
  wire [1:0] n2236_o;
  wire n2238_o;
  wire n2239_o;
  wire n2240_o;
  wire [1:0] n2241_o;
  wire n2243_o;
  wire [2:0] n2244_o;
  wire n2246_o;
  wire n2247_o;
  wire [1:0] n2248_o;
  wire n2250_o;
  wire n2251_o;
  wire n2252_o;
  wire [1:0] n2255_o;
  wire n2257_o;
  wire [1:0] n2258_o;
  wire n2260_o;
  wire n2263_o;
  wire n2266_o;
  wire n2268_o;
  wire [1:0] n2269_o;
  wire n2271_o;
  wire [1:0] n2274_o;
  wire n2275_o;
  wire n2276_o;
  wire n2279_o;
  wire n2280_o;
  wire n2281_o;
  wire n2282_o;
  wire [6:0] n2284_o;
  wire n2287_o;
  wire n2289_o;
  wire n2291_o;
  wire n2292_o;
  wire [1:0] n2293_o;
  wire n2295_o;
  wire n2298_o;
  wire n2301_o;
  wire n2303_o;
  wire n2305_o;
  wire n2307_o;
  wire n2309_o;
  wire n2311_o;
  wire n2313_o;
  wire n2314_o;
  wire [2:0] n2315_o;
  wire n2317_o;
  wire n2318_o;
  wire n2319_o;
  wire [1:0] n2320_o;
  wire n2322_o;
  wire [1:0] n2323_o;
  wire n2325_o;
  wire n2326_o;
  wire [2:0] n2327_o;
  wire n2329_o;
  wire [1:0] n2330_o;
  wire n2332_o;
  wire n2333_o;
  wire n2334_o;
  wire n2335_o;
  wire [5:0] n2336_o;
  wire n2338_o;
  wire n2339_o;
  wire n2340_o;
  wire [1:0] n2341_o;
  wire n2343_o;
  wire n2345_o;
  wire [1:0] n2346_o;
  reg [1:0] n2350_o;
  wire n2351_o;
  wire [5:0] n2352_o;
  wire n2354_o;
  wire n2355_o;
  wire n2357_o;
  wire n2358_o;
  wire [6:0] n2360_o;
  wire n2363_o;
  wire n2364_o;
  wire n2365_o;
  wire n2366_o;
  wire [6:0] n2368_o;
  wire n2370_o;
  wire n2371_o;
  wire [1:0] n2377_o;
  wire n2380_o;
  wire n2381_o;
  wire n2382_o;
  wire n2383_o;
  wire n2384_o;
  wire n2385_o;
  wire n2386_o;
  wire n2387_o;
  wire n2388_o;
  wire [6:0] n2390_o;
  wire [1:0] n2391_o;
  wire n2393_o;
  wire n2394_o;
  wire n2395_o;
  wire n2396_o;
  wire n2397_o;
  wire n2398_o;
  wire n2399_o;
  wire n2400_o;
  wire n2401_o;
  wire n2402_o;
  wire n2403_o;
  wire n2404_o;
  wire [6:0] n2405_o;
  wire [1:0] n2406_o;
  wire [1:0] n2407_o;
  wire n2409_o;
  wire n2412_o;
  wire n2415_o;
  wire n2416_o;
  wire n2417_o;
  wire n2418_o;
  wire n2419_o;
  wire n2420_o;
  wire n2421_o;
  wire n2422_o;
  wire n2423_o;
  wire n2424_o;
  wire n2425_o;
  wire n2426_o;
  wire n2427_o;
  wire [6:0] n2428_o;
  wire [1:0] n2429_o;
  wire n2431_o;
  wire [1:0] n2432_o;
  wire n2434_o;
  wire n2435_o;
  wire [2:0] n2436_o;
  wire n2438_o;
  wire n2439_o;
  wire [2:0] n2440_o;
  wire n2442_o;
  wire n2443_o;
  wire [3:0] n2444_o;
  wire n2446_o;
  wire n2447_o;
  wire [1:0] n2449_o;
  wire n2452_o;
  wire n2453_o;
  wire n2454_o;
  wire n2455_o;
  wire [6:0] n2457_o;
  wire n2458_o;
  wire n2461_o;
  wire n2462_o;
  wire n2463_o;
  wire n2464_o;
  wire n2466_o;
  wire n2467_o;
  wire n2470_o;
  wire n2473_o;
  wire [1:0] n2475_o;
  wire n2477_o;
  wire n2478_o;
  wire n2479_o;
  wire [6:0] n2481_o;
  wire [1:0] n2482_o;
  wire n2483_o;
  wire n2486_o;
  wire n2489_o;
  wire n2491_o;
  wire [1:0] n2492_o;
  wire n2494_o;
  wire [1:0] n2495_o;
  wire [1:0] n2496_o;
  wire n2498_o;
  wire n2500_o;
  wire n2502_o;
  wire [6:0] n2503_o;
  wire [1:0] n2504_o;
  wire [1:0] n2505_o;
  wire n2507_o;
  wire n2508_o;
  wire n2509_o;
  wire n2511_o;
  wire n2513_o;
  wire n2514_o;
  wire n2515_o;
  wire n2516_o;
  wire n2517_o;
  wire n2518_o;
  wire n2519_o;
  wire n2520_o;
  wire n2521_o;
  wire n2522_o;
  wire n2524_o;
  wire n2525_o;
  wire n2526_o;
  wire n2527_o;
  wire n2529_o;
  wire n2531_o;
  wire [6:0] n2532_o;
  wire [1:0] n2533_o;
  wire [1:0] n2534_o;
  wire n2536_o;
  wire n2538_o;
  wire n2540_o;
  wire n2542_o;
  wire [1:0] n2543_o;
  wire [1:0] n2544_o;
  wire n2546_o;
  wire n2547_o;
  wire n2548_o;
  wire [1:0] n2549_o;
  wire [1:0] n2550_o;
  wire [1:0] n2551_o;
  wire [1:0] n2552_o;
  wire n2553_o;
  wire n2554_o;
  wire n2555_o;
  wire n2556_o;
  wire n2558_o;
  wire n2560_o;
  wire [6:0] n2561_o;
  wire [2:0] n2562_o;
  wire n2564_o;
  wire n2565_o;
  wire [1:0] n2566_o;
  wire n2568_o;
  wire n2569_o;
  wire [1:0] n2570_o;
  wire n2572_o;
  wire n2573_o;
  wire [2:0] n2574_o;
  wire n2576_o;
  wire [1:0] n2577_o;
  wire n2579_o;
  wire n2580_o;
  wire n2581_o;
  wire n2584_o;
  wire n2587_o;
  wire n2589_o;
  wire n2591_o;
  wire [1:0] n2592_o;
  wire n2594_o;
  wire [2:0] n2595_o;
  wire n2597_o;
  wire n2598_o;
  wire [2:0] n2599_o;
  wire n2601_o;
  wire [2:0] n2602_o;
  wire n2604_o;
  wire [1:0] n2605_o;
  wire n2607_o;
  wire n2608_o;
  wire [2:0] n2609_o;
  wire n2611_o;
  wire n2612_o;
  wire n2613_o;
  wire n2614_o;
  wire n2615_o;
  wire n2619_o;
  wire n2622_o;
  wire n2624_o;
  wire n2626_o;
  wire n2628_o;
  wire n2630_o;
  wire [2:0] n2631_o;
  wire n2633_o;
  wire [2:0] n2634_o;
  wire n2636_o;
  wire [1:0] n2637_o;
  wire n2639_o;
  wire n2640_o;
  wire [2:0] n2641_o;
  wire n2643_o;
  wire n2644_o;
  wire n2645_o;
  wire n2646_o;
  wire n2647_o;
  wire n2650_o;
  wire n2652_o;
  wire n2654_o;
  wire n2655_o;
  wire n2656_o;
  wire n2658_o;
  wire [2:0] n2659_o;
  wire n2661_o;
  wire [2:0] n2662_o;
  wire n2664_o;
  wire n2665_o;
  wire [2:0] n2666_o;
  wire n2668_o;
  wire [1:0] n2669_o;
  wire n2671_o;
  wire n2672_o;
  wire n2675_o;
  wire n2677_o;
  wire n2679_o;
  wire n2680_o;
  wire n2681_o;
  wire n2683_o;
  wire [2:0] n2684_o;
  wire n2686_o;
  wire [2:0] n2687_o;
  wire n2689_o;
  wire [1:0] n2690_o;
  wire n2692_o;
  wire n2693_o;
  wire [2:0] n2694_o;
  wire n2696_o;
  wire n2697_o;
  wire n2698_o;
  wire n2699_o;
  wire n2700_o;
  wire n2703_o;
  wire n2705_o;
  wire n2707_o;
  wire n2708_o;
  wire n2709_o;
  wire n2711_o;
  wire [2:0] n2712_o;
  wire n2714_o;
  wire [2:0] n2715_o;
  wire n2717_o;
  wire n2718_o;
  wire n2719_o;
  wire n2720_o;
  wire n2723_o;
  wire n2725_o;
  wire n2727_o;
  wire n2728_o;
  wire n2729_o;
  wire n2731_o;
  wire n2732_o;
  wire n2733_o;
  wire n2734_o;
  wire n2735_o;
  wire n2736_o;
  wire n2737_o;
  wire n2738_o;
  wire n2739_o;
  wire n2740_o;
  wire n2741_o;
  wire n2742_o;
  wire [5:0] n2743_o;
  wire n2745_o;
  wire n2746_o;
  wire n2747_o;
  wire n2748_o;
  wire n2749_o;
  wire n2750_o;
  wire n2751_o;
  wire n2752_o;
  wire n2753_o;
  wire n2754_o;
  wire n2755_o;
  wire n2756_o;
  wire n2758_o;
  wire n2760_o;
  wire n2761_o;
  wire n2763_o;
  wire n2764_o;
  wire n2765_o;
  wire [1:0] n2767_o;
  wire [2:0] n2768_o;
  wire [1:0] n2769_o;
  wire [2:0] n2770_o;
  wire [2:0] n2771_o;
  wire [1:0] n2772_o;
  wire [1:0] n2773_o;
  wire [6:0] n2775_o;
  wire [1:0] n2776_o;
  wire n2779_o;
  wire n2781_o;
  wire [2:0] n2782_o;
  wire [2:0] n2783_o;
  wire n2784_o;
  wire n2785_o;
  wire [1:0] n2786_o;
  wire [1:0] n2787_o;
  wire [6:0] n2788_o;
  wire n2789_o;
  wire n2790_o;
  wire [5:0] n2791_o;
  wire n2793_o;
  wire n2794_o;
  wire n2795_o;
  wire n2796_o;
  wire n2797_o;
  wire n2798_o;
  wire n2799_o;
  wire n2800_o;
  wire n2801_o;
  wire n2805_o;
  wire n2807_o;
  wire n2809_o;
  wire n2810_o;
  wire n2811_o;
  wire n2812_o;
  wire n2813_o;
  wire n2814_o;
  wire [6:0] n2816_o;
  wire [1:0] n2817_o;
  wire n2819_o;
  wire n2822_o;
  wire [2:0] n2823_o;
  wire n2825_o;
  wire [1:0] n2826_o;
  wire n2828_o;
  wire n2831_o;
  wire n2834_o;
  wire n2836_o;
  wire [1:0] n2837_o;
  wire n2839_o;
  wire n2841_o;
  wire n2842_o;
  wire n2844_o;
  wire n2845_o;
  wire n2847_o;
  wire n2849_o;
  wire n2851_o;
  wire n2853_o;
  wire n2855_o;
  wire n2856_o;
  wire n2858_o;
  wire n2860_o;
  wire n2861_o;
  wire [1:0] n2862_o;
  wire n2864_o;
  wire n2865_o;
  wire n2866_o;
  wire n2868_o;
  wire n2869_o;
  wire [2:0] n2870_o;
  wire [2:0] n2871_o;
  wire n2872_o;
  wire n2873_o;
  wire n2874_o;
  wire n2875_o;
  wire [1:0] n2876_o;
  wire [1:0] n2877_o;
  wire n2878_o;
  wire n2879_o;
  wire n2880_o;
  wire n2881_o;
  wire n2882_o;
  wire n2884_o;
  wire n2886_o;
  wire [6:0] n2887_o;
  wire n2888_o;
  wire n2890_o;
  wire n2891_o;
  wire n2893_o;
  wire n2895_o;
  wire n2897_o;
  wire n2899_o;
  wire n2900_o;
  wire n2901_o;
  wire n2903_o;
  wire n2905_o;
  wire n2906_o;
  wire n2907_o;
  wire n2908_o;
  wire n2909_o;
  wire n2910_o;
  wire n2912_o;
  wire n2914_o;
  wire [6:0] n2915_o;
  wire n2916_o;
  wire n2918_o;
  wire n2919_o;
  wire n2921_o;
  wire n2923_o;
  wire n2925_o;
  wire n2927_o;
  wire n2929_o;
  wire n2931_o;
  wire n2933_o;
  wire n2935_o;
  wire n2937_o;
  wire n2938_o;
  wire [3:0] n2939_o;
  wire n2941_o;
  wire [3:0] n2943_o;
  wire n2945_o;
  wire n2947_o;
  wire n2948_o;
  wire [1:0] n2949_o;
  wire n2951_o;
  wire n2952_o;
  wire n2953_o;
  wire n2954_o;
  wire n2956_o;
  wire [2:0] n2957_o;
  wire [2:0] n2958_o;
  wire n2959_o;
  wire n2960_o;
  wire n2961_o;
  wire n2962_o;
  wire [1:0] n2963_o;
  wire [1:0] n2964_o;
  wire n2965_o;
  wire n2966_o;
  wire n2967_o;
  wire n2968_o;
  wire n2969_o;
  wire n2971_o;
  wire [3:0] n2973_o;
  wire n2975_o;
  wire n2977_o;
  wire [6:0] n2978_o;
  wire n2979_o;
  wire [1:0] n2980_o;
  wire n2982_o;
  wire n2984_o;
  wire n2985_o;
  wire n2986_o;
  wire n2988_o;
  wire n2989_o;
  wire n2991_o;
  wire [2:0] n2992_o;
  wire [2:0] n2993_o;
  wire n2995_o;
  wire n2997_o;
  wire n2998_o;
  wire n2999_o;
  wire n3000_o;
  wire n3001_o;
  wire n3002_o;
  wire n3003_o;
  wire n3004_o;
  wire [1:0] n3005_o;
  wire [1:0] n3006_o;
  wire n3007_o;
  wire n3008_o;
  wire n3009_o;
  wire n3010_o;
  wire n3011_o;
  wire n3012_o;
  wire n3013_o;
  wire n3015_o;
  wire n3017_o;
  wire n3019_o;
  wire n3021_o;
  wire [3:0] n3023_o;
  wire n3025_o;
  wire n3027_o;
  wire [6:0] n3028_o;
  wire [1:0] n3029_o;
  wire [1:0] n3030_o;
  wire n3031_o;
  wire n3033_o;
  wire n3034_o;
  wire n3035_o;
  wire n3037_o;
  wire n3038_o;
  wire n3040_o;
  wire n3042_o;
  wire [1:0] n3043_o;
  wire [1:0] n3044_o;
  wire [2:0] n3045_o;
  wire [2:0] n3046_o;
  wire n3047_o;
  wire n3048_o;
  wire n3049_o;
  wire n3050_o;
  wire n3051_o;
  wire n3052_o;
  wire n3053_o;
  wire n3054_o;
  wire n3055_o;
  wire n3056_o;
  wire n3057_o;
  wire [1:0] n3058_o;
  wire [1:0] n3059_o;
  wire [1:0] n3060_o;
  wire [1:0] n3061_o;
  wire n3062_o;
  wire n3063_o;
  wire n3064_o;
  wire n3065_o;
  wire n3066_o;
  wire n3067_o;
  wire n3068_o;
  wire n3069_o;
  wire n3071_o;
  wire [3:0] n3073_o;
  wire n3075_o;
  wire n3076_o;
  wire n3077_o;
  wire [6:0] n3078_o;
  wire [1:0] n3080_o;
  wire [1:0] n3081_o;
  wire n3083_o;
  wire n3085_o;
  wire n3087_o;
  wire n3088_o;
  wire n3090_o;
  wire n3092_o;
  wire n3094_o;
  wire n3096_o;
  wire n3098_o;
  wire [1:0] n3099_o;
  wire [1:0] n3100_o;
  wire [2:0] n3101_o;
  wire [2:0] n3102_o;
  wire n3103_o;
  wire n3104_o;
  wire n3105_o;
  wire n3106_o;
  wire n3107_o;
  wire n3108_o;
  wire [1:0] n3109_o;
  wire [1:0] n3110_o;
  wire n3111_o;
  wire n3112_o;
  wire n3113_o;
  wire n3114_o;
  wire [1:0] n3115_o;
  wire [1:0] n3116_o;
  wire [1:0] n3117_o;
  wire [1:0] n3118_o;
  wire n3119_o;
  wire n3120_o;
  wire n3121_o;
  wire n3122_o;
  wire n3123_o;
  wire n3124_o;
  wire n3125_o;
  wire n3126_o;
  wire n3127_o;
  wire n3129_o;
  wire n3131_o;
  wire [3:0] n3133_o;
  wire n3135_o;
  wire n3137_o;
  wire n3138_o;
  wire [6:0] n3139_o;
  wire n3141_o;
  wire [1:0] n3142_o;
  wire n3144_o;
  wire [2:0] n3145_o;
  wire n3147_o;
  wire n3148_o;
  wire [3:0] n3149_o;
  wire n3151_o;
  wire [1:0] n3152_o;
  wire n3154_o;
  wire n3155_o;
  wire n3156_o;
  wire n3157_o;
  wire [2:0] n3158_o;
  wire n3160_o;
  wire [2:0] n3161_o;
  wire n3163_o;
  wire n3164_o;
  wire n3165_o;
  wire n3166_o;
  wire [2:0] n3168_o;
  wire n3170_o;
  wire n3172_o;
  wire n3173_o;
  wire [1:0] n3174_o;
  wire n3176_o;
  wire [1:0] n3177_o;
  wire n3179_o;
  wire n3182_o;
  wire n3184_o;
  wire [1:0] n3185_o;
  wire n3187_o;
  wire n3189_o;
  wire [1:0] n3190_o;
  reg [1:0] n3194_o;
  wire n3195_o;
  wire n3198_o;
  wire [1:0] n3199_o;
  wire n3201_o;
  wire n3202_o;
  wire [2:0] n3203_o;
  wire n3205_o;
  wire n3208_o;
  wire n3210_o;
  wire n3213_o;
  wire n3215_o;
  wire [1:0] n3216_o;
  wire n3218_o;
  wire n3219_o;
  wire n3220_o;
  wire n3221_o;
  wire [2:0] n3222_o;
  wire n3225_o;
  wire n3227_o;
  wire n3228_o;
  wire n3229_o;
  wire [2:0] n3231_o;
  wire n3233_o;
  wire n3235_o;
  wire n3236_o;
  wire n3237_o;
  wire n3238_o;
  wire n3239_o;
  wire n3240_o;
  wire n3241_o;
  wire [2:0] n3243_o;
  wire n3245_o;
  wire n3247_o;
  wire n3248_o;
  wire n3249_o;
  wire n3250_o;
  wire n3251_o;
  wire n3252_o;
  wire n3253_o;
  wire n3255_o;
  wire n3256_o;
  wire n3258_o;
  wire n3260_o;
  wire n3261_o;
  wire n3263_o;
  wire n3264_o;
  wire n3266_o;
  wire n3268_o;
  wire [2:0] n3269_o;
  wire n3271_o;
  wire n3274_o;
  wire [1:0] n3275_o;
  reg n3276_o;
  reg [6:0] n3279_o;
  wire n3281_o;
  wire [4:0] n3282_o;
  reg [1:0] n3284_o;
  reg n3286_o;
  wire n3287_o;
  reg n3288_o;
  wire n3289_o;
  wire n3290_o;
  wire n3291_o;
  reg n3292_o;
  wire n3293_o;
  wire n3294_o;
  wire n3295_o;
  reg n3296_o;
  reg n3297_o;
  reg n3298_o;
  reg n3299_o;
  reg [6:0] n3303_o;
  wire [1:0] n3304_o;
  wire n3305_o;
  wire [1:0] n3306_o;
  wire n3307_o;
  wire n3308_o;
  wire [1:0] n3309_o;
  wire n3310_o;
  wire n3311_o;
  wire n3312_o;
  wire [6:0] n3313_o;
  wire [1:0] n3314_o;
  wire n3315_o;
  wire n3316_o;
  wire n3318_o;
  wire n3321_o;
  wire n3323_o;
  wire n3325_o;
  wire n3328_o;
  wire n3331_o;
  wire n3334_o;
  wire [1:0] n3335_o;
  wire n3337_o;
  wire n3338_o;
  wire n3339_o;
  wire [1:0] n3340_o;
  wire [1:0] n3341_o;
  wire n3342_o;
  wire n3344_o;
  wire n3346_o;
  wire n3347_o;
  wire n3349_o;
  wire n3351_o;
  wire n3352_o;
  wire n3354_o;
  wire n3355_o;
  wire n3356_o;
  wire n3357_o;
  wire [2:0] n3358_o;
  wire n3360_o;
  wire [2:0] n3361_o;
  wire n3363_o;
  wire n3364_o;
  wire n3365_o;
  wire n3366_o;
  wire n3367_o;
  wire n3374_o;
  wire n3377_o;
  wire n3380_o;
  wire n3382_o;
  wire n3384_o;
  wire n3386_o;
  wire n3388_o;
  wire n3389_o;
  wire n3390_o;
  wire [1:0] n3391_o;
  wire n3393_o;
  wire n3394_o;
  wire n3395_o;
  wire [2:0] n3396_o;
  wire n3398_o;
  wire n3399_o;
  wire [3:0] n3400_o;
  wire n3402_o;
  wire n3403_o;
  wire [2:0] n3407_o;
  wire n3409_o;
  wire n3412_o;
  wire n3415_o;
  wire n3418_o;
  wire n3419_o;
  wire [1:0] n3421_o;
  wire n3423_o;
  wire n3425_o;
  wire n3427_o;
  wire n3428_o;
  wire n3431_o;
  wire n3434_o;
  wire n3437_o;
  wire n3439_o;
  wire n3441_o;
  wire n3442_o;
  wire n3445_o;
  wire n3448_o;
  wire n3450_o;
  wire n3451_o;
  wire n3452_o;
  wire n3454_o;
  wire n3456_o;
  wire [1:0] n3457_o;
  wire n3459_o;
  wire n3461_o;
  wire n3462_o;
  wire n3464_o;
  wire n3466_o;
  wire n3467_o;
  wire n3468_o;
  wire n3469_o;
  wire n3471_o;
  wire n3472_o;
  wire n3473_o;
  wire n3474_o;
  wire n3476_o;
  wire n3477_o;
  wire n3479_o;
  wire [2:0] n3480_o;
  wire n3482_o;
  wire [3:0] n3483_o;
  wire n3485_o;
  wire [1:0] n3486_o;
  wire n3488_o;
  wire n3489_o;
  wire n3490_o;
  wire n3491_o;
  wire n3493_o;
  wire n3494_o;
  wire n3495_o;
  wire n3496_o;
  wire n3497_o;
  wire n3498_o;
  wire n3499_o;
  wire n3500_o;
  wire n3503_o;
  wire n3504_o;
  wire n3506_o;
  wire n3507_o;
  wire n3508_o;
  wire n3509_o;
  wire n3510_o;
  wire n3511_o;
  wire n3512_o;
  wire n3513_o;
  wire n3516_o;
  wire [1:0] n3518_o;
  wire n3521_o;
  wire n3523_o;
  wire n3524_o;
  wire n3525_o;
  wire [1:0] n3527_o;
  wire n3529_o;
  wire n3530_o;
  wire n3531_o;
  wire n3532_o;
  wire n3533_o;
  wire n3534_o;
  wire [1:0] n3535_o;
  wire n3537_o;
  wire n3538_o;
  wire n3539_o;
  wire n3540_o;
  wire n3541_o;
  wire n3543_o;
  wire n3544_o;
  wire n3547_o;
  wire n3551_o;
  wire n3554_o;
  wire n3556_o;
  wire n3558_o;
  wire n3561_o;
  wire n3562_o;
  wire n3563_o;
  wire n3565_o;
  wire [1:0] n3566_o;
  wire n3568_o;
  wire n3570_o;
  wire n3572_o;
  wire n3574_o;
  wire n3576_o;
  wire n3577_o;
  wire n3578_o;
  wire n3580_o;
  wire n3582_o;
  wire [1:0] n3583_o;
  wire [1:0] n3584_o;
  wire n3586_o;
  wire n3588_o;
  wire n3589_o;
  wire n3591_o;
  wire n3592_o;
  wire n3593_o;
  wire n3594_o;
  wire n3595_o;
  wire n3596_o;
  wire n3597_o;
  wire n3598_o;
  wire n3599_o;
  wire n3600_o;
  wire n3601_o;
  wire n3602_o;
  wire n3604_o;
  wire n3606_o;
  wire n3608_o;
  wire n3610_o;
  wire n3612_o;
  wire [2:0] n3613_o;
  wire [2:0] n3614_o;
  wire n3616_o;
  wire [2:0] n3617_o;
  wire n3619_o;
  wire [1:0] n3620_o;
  wire n3622_o;
  wire n3623_o;
  wire n3624_o;
  wire [1:0] n3625_o;
  wire n3627_o;
  wire n3629_o;
  wire n3631_o;
  wire n3632_o;
  wire n3633_o;
  wire n3634_o;
  wire n3636_o;
  wire [1:0] n3637_o;
  wire n3639_o;
  wire n3642_o;
  wire [1:0] n3646_o;
  wire n3648_o;
  wire n3651_o;
  wire n3653_o;
  wire n3654_o;
  wire n3655_o;
  wire [1:0] n3657_o;
  wire n3660_o;
  wire n3661_o;
  wire n3662_o;
  wire n3663_o;
  wire n3664_o;
  wire n3666_o;
  wire n3668_o;
  wire n3670_o;
  wire n3671_o;
  wire n3672_o;
  wire n3673_o;
  wire n3676_o;
  wire n3678_o;
  wire n3681_o;
  wire n3684_o;
  wire n3687_o;
  wire n3688_o;
  wire n3689_o;
  wire n3690_o;
  wire n3691_o;
  wire [1:0] n3692_o;
  wire [1:0] n3694_o;
  wire n3696_o;
  wire n3698_o;
  wire n3700_o;
  wire [2:0] n3701_o;
  wire n3703_o;
  wire [2:0] n3704_o;
  wire n3706_o;
  wire [1:0] n3707_o;
  wire n3709_o;
  wire n3710_o;
  wire n3711_o;
  wire [1:0] n3712_o;
  wire n3714_o;
  wire n3717_o;
  wire n3719_o;
  wire n3720_o;
  wire n3721_o;
  wire n3722_o;
  wire n3724_o;
  wire n3726_o;
  wire n3727_o;
  wire [1:0] n3728_o;
  wire n3730_o;
  wire n3733_o;
  wire n3734_o;
  wire n3737_o;
  wire n3740_o;
  wire n3743_o;
  wire n3746_o;
  wire n3747_o;
  wire n3748_o;
  wire n3750_o;
  wire n3752_o;
  wire n3753_o;
  wire n3755_o;
  wire n3757_o;
  wire n3759_o;
  wire n3761_o;
  wire n3762_o;
  wire n3763_o;
  wire n3765_o;
  wire n3767_o;
  wire n3769_o;
  wire [1:0] n3770_o;
  wire n3772_o;
  wire [2:0] n3773_o;
  wire n3775_o;
  wire [3:0] n3776_o;
  wire n3778_o;
  wire [1:0] n3779_o;
  wire n3781_o;
  wire n3782_o;
  wire n3783_o;
  wire [1:0] n3784_o;
  wire n3786_o;
  wire n3787_o;
  wire n3789_o;
  wire n3790_o;
  wire n3791_o;
  wire n3792_o;
  wire n3793_o;
  wire n3795_o;
  wire n3796_o;
  wire [1:0] n3798_o;
  wire n3801_o;
  wire n3804_o;
  wire n3807_o;
  wire n3810_o;
  wire n3812_o;
  wire [2:0] n3813_o;
  wire n3815_o;
  wire [2:0] n3816_o;
  wire n3818_o;
  wire [1:0] n3819_o;
  wire n3821_o;
  wire n3822_o;
  wire n3823_o;
  wire [1:0] n3826_o;
  wire n3828_o;
  wire n3831_o;
  wire n3833_o;
  wire n3834_o;
  wire n3837_o;
  wire n3840_o;
  wire n3843_o;
  wire n3846_o;
  wire n3849_o;
  wire n3851_o;
  wire n3852_o;
  wire n3853_o;
  wire n3855_o;
  wire n3857_o;
  wire n3858_o;
  wire n3860_o;
  wire n3861_o;
  wire n3862_o;
  wire n3863_o;
  wire n3864_o;
  wire n3866_o;
  wire n3867_o;
  wire n3868_o;
  wire n3869_o;
  wire n3870_o;
  wire n3872_o;
  wire n3874_o;
  wire n3876_o;
  wire [1:0] n3877_o;
  wire n3879_o;
  wire [2:0] n3880_o;
  wire n3882_o;
  wire [3:0] n3883_o;
  wire n3885_o;
  wire [1:0] n3886_o;
  wire n3888_o;
  wire n3889_o;
  wire n3890_o;
  wire [1:0] n3891_o;
  wire n3893_o;
  wire n3894_o;
  wire n3896_o;
  wire n3897_o;
  wire n3898_o;
  wire n3899_o;
  wire n3900_o;
  wire [1:0] n3903_o;
  wire [1:0] n3904_o;
  wire [1:0] n3905_o;
  wire n3906_o;
  wire [1:0] n3907_o;
  wire n3909_o;
  wire n3910_o;
  wire n3911_o;
  wire n3913_o;
  wire n3914_o;
  wire n3915_o;
  wire n3916_o;
  wire n3917_o;
  wire [1:0] n3919_o;
  wire [1:0] n3921_o;
  wire n3922_o;
  wire n3925_o;
  wire n3928_o;
  wire n3931_o;
  wire n3934_o;
  wire n3936_o;
  wire n3937_o;
  wire n3938_o;
  wire n3940_o;
  wire n3943_o;
  wire n3945_o;
  wire n3947_o;
  wire n3949_o;
  wire n3951_o;
  wire [2:0] n3952_o;
  wire n3954_o;
  wire [2:0] n3955_o;
  wire n3957_o;
  wire [1:0] n3958_o;
  wire n3960_o;
  wire n3961_o;
  wire n3962_o;
  wire [2:0] n3965_o;
  wire n3967_o;
  wire n3970_o;
  wire n3972_o;
  wire n3973_o;
  wire n3976_o;
  wire n3979_o;
  wire n3982_o;
  wire n3985_o;
  wire n3987_o;
  wire n3989_o;
  wire n3991_o;
  wire n3993_o;
  wire n3994_o;
  wire n3995_o;
  wire n3997_o;
  wire n3999_o;
  wire n4000_o;
  wire n4002_o;
  wire n4003_o;
  wire n4004_o;
  wire n4006_o;
  wire n4007_o;
  wire n4008_o;
  wire n4010_o;
  wire n4012_o;
  wire n4014_o;
  wire n4016_o;
  wire n4017_o;
  wire [2:0] n4018_o;
  wire n4020_o;
  wire n4021_o;
  wire n4022_o;
  wire n4023_o;
  wire n4027_o;
  wire n4028_o;
  wire [1:0] n4031_o;
  wire n4033_o;
  wire n4034_o;
  wire n4035_o;
  wire [1:0] n4036_o;
  wire n4038_o;
  wire n4039_o;
  wire [2:0] n4040_o;
  wire n4042_o;
  wire [1:0] n4043_o;
  wire n4045_o;
  wire n4046_o;
  wire n4047_o;
  wire n4048_o;
  wire n4049_o;
  wire n4050_o;
  wire [1:0] n4051_o;
  wire n4053_o;
  wire [2:0] n4054_o;
  wire n4056_o;
  wire n4057_o;
  wire [3:0] n4058_o;
  wire n4060_o;
  wire n4061_o;
  wire n4062_o;
  wire n4063_o;
  wire n4065_o;
  wire n4066_o;
  wire [1:0] n4068_o;
  wire [2:0] n4069_o;
  wire n4071_o;
  wire [2:0] n4072_o;
  wire n4074_o;
  wire n4075_o;
  wire n4077_o;
  wire n4078_o;
  wire n4082_o;
  wire n4084_o;
  wire [2:0] n4085_o;
  wire n4087_o;
  wire n4091_o;
  wire n4092_o;
  wire n4093_o;
  wire n4095_o;
  wire n4096_o;
  wire n4097_o;
  wire n4100_o;
  wire n4101_o;
  wire n4102_o;
  wire n4103_o;
  wire [2:0] n4105_o;
  wire n4107_o;
  wire [2:0] n4108_o;
  wire n4110_o;
  wire n4111_o;
  wire [2:0] n4112_o;
  wire n4114_o;
  wire n4115_o;
  wire n4117_o;
  wire n4118_o;
  wire [6:0] n4121_o;
  wire n4122_o;
  wire n4123_o;
  wire n4124_o;
  wire n4125_o;
  wire [6:0] n4126_o;
  wire n4127_o;
  wire n4129_o;
  wire n4130_o;
  wire [1:0] n4134_o;
  wire n4135_o;
  wire n4136_o;
  wire [1:0] n4139_o;
  wire n4141_o;
  wire n4142_o;
  wire n4143_o;
  wire n4144_o;
  wire n4145_o;
  wire [6:0] n4147_o;
  wire [1:0] n4148_o;
  wire n4150_o;
  wire n4152_o;
  wire n4154_o;
  wire n4155_o;
  wire n4156_o;
  wire n4157_o;
  wire n4160_o;
  wire n4162_o;
  wire n4165_o;
  wire n4168_o;
  wire [1:0] n4169_o;
  wire n4171_o;
  wire n4173_o;
  wire n4175_o;
  wire n4177_o;
  wire [1:0] n4178_o;
  wire n4180_o;
  wire n4182_o;
  wire n4184_o;
  wire n4186_o;
  wire n4188_o;
  wire [6:0] n4189_o;
  wire [1:0] n4190_o;
  wire [1:0] n4191_o;
  wire n4193_o;
  wire n4196_o;
  wire n4198_o;
  wire n4200_o;
  wire n4202_o;
  wire n4203_o;
  wire n4204_o;
  wire n4205_o;
  wire n4206_o;
  wire n4207_o;
  wire n4208_o;
  wire n4209_o;
  wire n4210_o;
  wire [1:0] n4211_o;
  wire n4212_o;
  wire n4213_o;
  wire n4214_o;
  wire n4215_o;
  wire n4216_o;
  wire n4217_o;
  wire n4219_o;
  wire n4221_o;
  wire n4223_o;
  wire n4224_o;
  wire n4226_o;
  wire [6:0] n4227_o;
  wire n4228_o;
  wire [1:0] n4244_o;
  wire n4246_o;
  wire [2:0] n4247_o;
  wire n4249_o;
  wire n4250_o;
  wire [3:0] n4251_o;
  wire n4253_o;
  wire [1:0] n4254_o;
  wire n4256_o;
  wire n4257_o;
  wire n4258_o;
  wire n4259_o;
  wire n4260_o;
  wire n4262_o;
  wire n4264_o;
  wire n4265_o;
  wire n4266_o;
  wire n4267_o;
  wire n4268_o;
  wire n4270_o;
  wire n4272_o;
  wire n4273_o;
  wire n4274_o;
  wire n4275_o;
  wire n4278_o;
  wire n4279_o;
  wire n4280_o;
  wire n4281_o;
  wire [6:0] n4283_o;
  wire n4285_o;
  wire n4286_o;
  wire [1:0] n4287_o;
  wire n4289_o;
  wire n4290_o;
  wire n4291_o;
  wire n4292_o;
  wire n4293_o;
  wire n4295_o;
  wire n4296_o;
  wire [6:0] n4299_o;
  wire [1:0] n4301_o;
  wire n4304_o;
  wire n4307_o;
  wire n4308_o;
  wire n4309_o;
  wire [6:0] n4310_o;
  wire [1:0] n4311_o;
  wire n4313_o;
  wire n4314_o;
  wire n4315_o;
  wire n4318_o;
  wire [1:0] n4320_o;
  wire n4321_o;
  wire n4324_o;
  wire n4326_o;
  wire n4328_o;
  wire n4330_o;
  wire n4333_o;
  wire n4336_o;
  wire n4338_o;
  wire n4340_o;
  wire n4342_o;
  wire [6:0] n4343_o;
  wire n4344_o;
  wire [2:0] n4345_o;
  wire n4347_o;
  wire [2:0] n4350_o;
  wire n4352_o;
  wire n4353_o;
  wire [1:0] n4354_o;
  wire n4356_o;
  wire n4357_o;
  wire [2:0] n4358_o;
  wire n4360_o;
  wire n4361_o;
  wire [3:0] n4362_o;
  wire n4364_o;
  wire n4365_o;
  wire n4367_o;
  wire n4368_o;
  wire [1:0] n4371_o;
  wire n4373_o;
  wire n4374_o;
  wire n4375_o;
  wire n4376_o;
  wire n4377_o;
  wire [6:0] n4379_o;
  wire n4380_o;
  wire [1:0] n4382_o;
  wire [1:0] n4383_o;
  wire n4384_o;
  wire n4387_o;
  wire n4390_o;
  wire n4393_o;
  wire n4396_o;
  wire n4397_o;
  wire n4398_o;
  wire n4399_o;
  wire n4400_o;
  wire n4401_o;
  wire [1:0] n4402_o;
  wire n4403_o;
  wire n4405_o;
  wire n4407_o;
  wire n4409_o;
  wire n4411_o;
  wire n4412_o;
  wire n4413_o;
  wire n4414_o;
  wire n4415_o;
  wire [6:0] n4416_o;
  wire [1:0] n4417_o;
  wire n4418_o;
  wire n4420_o;
  wire n4422_o;
  wire n4424_o;
  wire n4426_o;
  wire n4427_o;
  wire n4428_o;
  wire n4429_o;
  wire n4430_o;
  wire n4432_o;
  wire n4434_o;
  wire [6:0] n4435_o;
  wire [2:0] n4436_o;
  wire n4438_o;
  wire n4448_o;
  wire n4451_o;
  wire n4454_o;
  wire n4455_o;
  wire n4456_o;
  wire n4457_o;
  wire n4458_o;
  wire n4459_o;
  wire n4460_o;
  wire n4461_o;
  wire n4462_o;
  wire n4463_o;
  wire n4464_o;
  wire n4465_o;
  wire [6:0] n4467_o;
  wire [2:0] n4468_o;
  wire n4470_o;
  wire [2:0] n4471_o;
  wire n4473_o;
  wire [1:0] n4474_o;
  wire n4476_o;
  wire n4477_o;
  wire n4478_o;
  wire [1:0] n4483_o;
  wire n4485_o;
  wire n4488_o;
  wire n4490_o;
  wire n4491_o;
  wire n4494_o;
  wire n4497_o;
  wire n4500_o;
  wire n4503_o;
  wire n4506_o;
  wire n4508_o;
  wire n4509_o;
  wire n4510_o;
  wire n4512_o;
  wire n4514_o;
  wire n4516_o;
  wire n4518_o;
  wire [1:0] n4520_o;
  wire n4522_o;
  wire n4523_o;
  wire n4525_o;
  wire n4526_o;
  wire n4528_o;
  wire n4530_o;
  wire n4532_o;
  wire n4534_o;
  wire n4536_o;
  wire n4537_o;
  wire n4538_o;
  wire n4539_o;
  wire n4540_o;
  wire n4541_o;
  wire n4542_o;
  wire n4543_o;
  wire n4544_o;
  wire n4546_o;
  wire n4547_o;
  wire n4548_o;
  wire n4549_o;
  wire n4550_o;
  wire n4552_o;
  wire n4554_o;
  wire n4555_o;
  wire n4556_o;
  wire [1:0] n4558_o;
  wire [1:0] n4559_o;
  wire n4561_o;
  wire n4562_o;
  wire n4564_o;
  wire n4566_o;
  wire n4568_o;
  wire n4569_o;
  wire n4570_o;
  wire n4571_o;
  wire [2:0] n4572_o;
  wire n4573_o;
  wire n4574_o;
  wire n4575_o;
  wire n4576_o;
  wire n4577_o;
  wire n4578_o;
  wire n4579_o;
  wire [2:0] n4580_o;
  wire [2:0] n4581_o;
  wire n4582_o;
  wire n4584_o;
  wire n4586_o;
  wire n4588_o;
  wire n4590_o;
  wire n4591_o;
  wire [6:0] n4592_o;
  wire [1:0] n4593_o;
  wire [1:0] n4594_o;
  wire n4596_o;
  wire n4597_o;
  wire n4599_o;
  wire n4601_o;
  wire n4602_o;
  wire n4604_o;
  wire n4606_o;
  wire n4608_o;
  wire n4609_o;
  wire n4610_o;
  wire n4612_o;
  wire n4614_o;
  wire n4615_o;
  wire n4616_o;
  wire n4618_o;
  wire n4619_o;
  wire n4620_o;
  wire n4621_o;
  wire n4622_o;
  wire n4623_o;
  wire n4624_o;
  wire n4625_o;
  wire n4626_o;
  wire [2:0] n4627_o;
  wire [2:0] n4628_o;
  wire n4630_o;
  wire n4631_o;
  wire n4633_o;
  wire n4635_o;
  wire n4637_o;
  wire n4639_o;
  wire n4641_o;
  wire [6:0] n4642_o;
  wire [1:0] n4643_o;
  wire [1:0] n4644_o;
  wire n4646_o;
  wire n4647_o;
  wire n4648_o;
  wire n4650_o;
  wire n4651_o;
  wire n4653_o;
  wire n4655_o;
  wire n4657_o;
  wire n4659_o;
  wire n4660_o;
  wire n4661_o;
  wire n4663_o;
  wire n4664_o;
  wire n4665_o;
  wire n4666_o;
  wire n4667_o;
  wire n4668_o;
  wire n4669_o;
  wire n4670_o;
  wire n4671_o;
  wire n4672_o;
  wire n4673_o;
  wire n4674_o;
  wire n4675_o;
  wire n4676_o;
  wire n4677_o;
  wire n4678_o;
  wire n4679_o;
  wire n4680_o;
  wire n4681_o;
  wire n4682_o;
  wire n4683_o;
  wire n4684_o;
  wire n4685_o;
  wire n4686_o;
  wire n4687_o;
  wire n4688_o;
  wire n4689_o;
  wire n4690_o;
  wire n4691_o;
  wire n4692_o;
  wire n4693_o;
  wire n4694_o;
  wire n4695_o;
  wire n4696_o;
  wire n4697_o;
  wire n4699_o;
  wire n4701_o;
  wire n4703_o;
  wire n4705_o;
  wire n4707_o;
  wire n4709_o;
  wire n4711_o;
  wire n4712_o;
  wire n4714_o;
  wire [6:0] n4715_o;
  wire n4717_o;
  wire n4719_o;
  wire n4720_o;
  wire [4:0] n4721_o;
  wire n4723_o;
  wire [1:0] n4724_o;
  wire n4726_o;
  wire n4727_o;
  wire [1:0] n4728_o;
  wire n4730_o;
  wire [2:0] n4731_o;
  wire n4733_o;
  wire [2:0] n4734_o;
  wire n4736_o;
  wire [1:0] n4737_o;
  wire n4739_o;
  wire n4740_o;
  wire n4741_o;
  wire n4742_o;
  wire [1:0] n4743_o;
  wire n4745_o;
  wire [2:0] n4746_o;
  wire n4748_o;
  wire n4749_o;
  wire [3:0] n4750_o;
  wire n4752_o;
  wire [1:0] n4753_o;
  wire n4755_o;
  wire n4756_o;
  wire n4757_o;
  wire n4758_o;
  wire n4759_o;
  wire n4762_o;
  wire n4764_o;
  wire n4767_o;
  wire [1:0] n4769_o;
  wire n4771_o;
  wire [1:0] n4772_o;
  wire n4774_o;
  wire n4777_o;
  wire [1:0] n4779_o;
  wire n4782_o;
  wire n4785_o;
  wire n4787_o;
  wire n4788_o;
  wire n4790_o;
  wire n4792_o;
  wire n4794_o;
  wire n4796_o;
  wire n4799_o;
  wire n4802_o;
  wire n4805_o;
  wire n4807_o;
  wire n4809_o;
  wire [1:0] n4810_o;
  wire n4812_o;
  wire n4814_o;
  wire n4816_o;
  wire n4818_o;
  wire n4820_o;
  wire n4822_o;
  wire n4824_o;
  wire n4826_o;
  wire n4828_o;
  wire n4830_o;
  wire n4831_o;
  wire n4832_o;
  wire [1:0] n4833_o;
  wire n4835_o;
  wire n4836_o;
  wire [2:0] n4837_o;
  wire n4839_o;
  wire n4840_o;
  wire [3:0] n4841_o;
  wire n4843_o;
  wire n4844_o;
  wire n4845_o;
  wire [6:0] n4847_o;
  wire n4849_o;
  wire n4850_o;
  wire n4851_o;
  wire n4852_o;
  wire n4853_o;
  wire [1:0] n4856_o;
  wire n4858_o;
  wire n4859_o;
  wire n4860_o;
  wire n4861_o;
  wire n4862_o;
  wire [6:0] n4864_o;
  wire n4866_o;
  wire n4867_o;
  wire n4868_o;
  wire n4869_o;
  wire n4871_o;
  wire n4873_o;
  wire n4876_o;
  wire n4878_o;
  wire n4879_o;
  wire n4880_o;
  wire n4881_o;
  wire n4883_o;
  wire n4885_o;
  wire [1:0] n4887_o;
  wire n4888_o;
  wire n4889_o;
  wire n4890_o;
  wire [1:0] n4892_o;
  wire [1:0] n4893_o;
  wire n4894_o;
  wire n4896_o;
  wire n4899_o;
  wire n4902_o;
  wire n4905_o;
  wire n4908_o;
  wire [1:0] n4909_o;
  wire n4910_o;
  wire n4911_o;
  wire n4912_o;
  wire n4913_o;
  wire [1:0] n4914_o;
  wire [6:0] n4915_o;
  wire [6:0] n4916_o;
  wire n4918_o;
  wire n4920_o;
  wire n4921_o;
  wire n4923_o;
  wire n4924_o;
  wire n4926_o;
  wire n4927_o;
  wire n4929_o;
  wire n4930_o;
  wire n4932_o;
  wire n4933_o;
  wire n4935_o;
  wire n4936_o;
  wire n4938_o;
  wire n4939_o;
  wire n4941_o;
  wire n4942_o;
  wire n4944_o;
  wire n4945_o;
  wire n4947_o;
  wire n4948_o;
  wire n4950_o;
  wire n4951_o;
  wire n4953_o;
  wire n4954_o;
  wire n4956_o;
  wire n4957_o;
  wire n4959_o;
  wire n4960_o;
  wire n4962_o;
  wire n4963_o;
  wire n4971_o;
  wire n4974_o;
  wire n4977_o;
  wire n4978_o;
  wire n4979_o;
  wire n4980_o;
  wire n4981_o;
  wire n4982_o;
  wire n4983_o;
  wire n4984_o;
  wire n4985_o;
  wire [6:0] n4987_o;
  wire n4989_o;
  wire n4991_o;
  wire n4992_o;
  wire n4994_o;
  wire n4995_o;
  wire n4997_o;
  wire n4998_o;
  wire n5000_o;
  wire n5001_o;
  wire n5003_o;
  wire n5004_o;
  wire n5006_o;
  wire n5007_o;
  wire n5009_o;
  wire n5010_o;
  wire [1:0] n5017_o;
  wire n5019_o;
  wire n5022_o;
  wire n5025_o;
  wire n5026_o;
  wire n5027_o;
  wire n5028_o;
  wire n5029_o;
  wire [6:0] n5031_o;
  wire n5033_o;
  wire n5035_o;
  wire n5036_o;
  wire n5038_o;
  wire n5039_o;
  wire n5041_o;
  wire n5042_o;
  wire n5044_o;
  wire n5045_o;
  wire n5047_o;
  wire n5048_o;
  wire n5050_o;
  wire n5051_o;
  wire n5053_o;
  wire n5054_o;
  wire [1:0] n5057_o;
  wire n5060_o;
  wire n5063_o;
  wire n5066_o;
  wire n5069_o;
  wire n5070_o;
  wire n5071_o;
  wire n5072_o;
  wire n5073_o;
  wire n5075_o;
  wire n5077_o;
  wire n5078_o;
  wire n5080_o;
  wire n5081_o;
  wire n5083_o;
  wire n5084_o;
  wire n5086_o;
  wire n5087_o;
  wire n5089_o;
  wire n5090_o;
  wire n5092_o;
  wire n5093_o;
  wire n5095_o;
  wire n5096_o;
  wire [1:0] n5100_o;
  wire n5103_o;
  wire n5106_o;
  wire n5107_o;
  wire n5108_o;
  wire n5109_o;
  wire n5110_o;
  wire n5112_o;
  wire n5114_o;
  wire n5116_o;
  wire n5117_o;
  wire n5119_o;
  wire n5120_o;
  wire n5122_o;
  wire n5123_o;
  wire n5125_o;
  wire n5126_o;
  wire n5128_o;
  wire n5129_o;
  wire n5131_o;
  wire n5132_o;
  wire n5134_o;
  wire n5135_o;
  wire n5136_o;
  wire [5:0] n5140_o;
  wire n5141_o;
  wire n5142_o;
  wire [5:0] n5143_o;
  wire n5146_o;
  wire n5149_o;
  wire n5150_o;
  wire n5151_o;
  wire n5152_o;
  wire n5153_o;
  wire n5155_o;
  wire n5157_o;
  wire n5158_o;
  wire n5160_o;
  wire n5163_o;
  wire n5165_o;
  wire n5166_o;
  wire n5167_o;
  wire n5170_o;
  wire n5173_o;
  wire n5175_o;
  wire n5177_o;
  wire n5178_o;
  wire n5179_o;
  wire n5181_o;
  wire n5184_o;
  wire n5185_o;
  wire n5186_o;
  wire n5187_o;
  wire [1:0] n5189_o;
  wire n5191_o;
  wire [1:0] n5192_o;
  wire n5193_o;
  wire n5194_o;
  wire n5195_o;
  wire n5196_o;
  wire [1:0] n5197_o;
  wire [1:0] n5198_o;
  wire [6:0] n5200_o;
  wire n5201_o;
  wire n5202_o;
  wire n5205_o;
  wire n5208_o;
  wire n5209_o;
  wire n5210_o;
  wire n5211_o;
  wire n5212_o;
  wire n5214_o;
  wire n5215_o;
  wire n5217_o;
  wire n5219_o;
  wire n5220_o;
  wire [1:0] n5225_o;
  wire n5227_o;
  wire n5229_o;
  wire [1:0] n5230_o;
  wire n5231_o;
  wire n5232_o;
  wire n5233_o;
  wire n5234_o;
  wire [1:0] n5235_o;
  wire [1:0] n5236_o;
  wire [6:0] n5238_o;
  wire n5240_o;
  wire [1:0] n5245_o;
  wire n5247_o;
  wire [1:0] n5248_o;
  wire n5249_o;
  wire n5250_o;
  wire n5251_o;
  wire n5252_o;
  wire [1:0] n5253_o;
  wire [1:0] n5254_o;
  wire [6:0] n5256_o;
  wire n5258_o;
  wire [1:0] n5260_o;
  wire n5261_o;
  wire n5263_o;
  wire n5264_o;
  wire n5267_o;
  wire n5270_o;
  wire n5272_o;
  wire n5274_o;
  wire n5275_o;
  wire [11:0] n5276_o;
  wire n5278_o;
  wire n5280_o;
  wire n5282_o;
  wire n5283_o;
  wire n5284_o;
  wire n5285_o;
  wire [1:0] n5286_o;
  wire [1:0] n5287_o;
  wire n5288_o;
  wire n5289_o;
  wire n5293_o;
  wire n5295_o;
  wire n5297_o;
  wire [6:0] n5299_o;
  wire [1:0] n5301_o;
  wire n5302_o;
  wire n5305_o;
  wire n5308_o;
  wire [1:0] n5309_o;
  wire [1:0] n5310_o;
  wire [1:0] n5312_o;
  wire [6:0] n5313_o;
  wire [1:0] n5314_o;
  wire n5315_o;
  wire n5318_o;
  wire n5320_o;
  wire n5322_o;
  wire [1:0] n5323_o;
  wire [1:0] n5325_o;
  wire [6:0] n5326_o;
  wire n5328_o;
  wire n5330_o;
  wire n5331_o;
  wire [12:0] n5332_o;
  reg n5333_o;
  reg [1:0] n5338_o;
  reg [1:0] n5339_o;
  reg n5340_o;
  reg n5341_o;
  reg n5342_o;
  reg n5344_o;
  reg n5346_o;
  reg [5:0] n5347_o;
  reg n5348_o;
  reg n5351_o;
  reg n5353_o;
  reg n5356_o;
  reg n5358_o;
  reg n5362_o;
  reg n5364_o;
  wire n5365_o;
  reg n5366_o;
  wire n5367_o;
  reg n5368_o;
  wire n5369_o;
  reg n5370_o;
  wire n5371_o;
  reg n5372_o;
  wire n5373_o;
  wire n5374_o;
  wire n5375_o;
  reg n5376_o;
  wire n5377_o;
  wire n5378_o;
  wire n5379_o;
  reg n5380_o;
  wire n5381_o;
  reg n5382_o;
  wire n5383_o;
  reg n5384_o;
  wire [1:0] n5385_o;
  reg [1:0] n5386_o;
  wire [1:0] n5387_o;
  reg [1:0] n5388_o;
  wire n5389_o;
  wire n5390_o;
  wire n5391_o;
  wire n5392_o;
  reg n5393_o;
  wire n5394_o;
  wire n5395_o;
  wire n5396_o;
  wire n5397_o;
  reg n5398_o;
  wire n5399_o;
  reg n5400_o;
  reg n5402_o;
  reg n5404_o;
  reg [1:0] n5406_o;
  reg n5408_o;
  reg [6:0] n5409_o;
  wire n5410_o;
  wire [1:0] n5411_o;
  wire [1:0] n5412_o;
  wire n5413_o;
  wire n5414_o;
  wire n5415_o;
  wire n5417_o;
  wire n5419_o;
  wire n5421_o;
  wire n5423_o;
  wire [5:0] n5424_o;
  wire n5425_o;
  wire n5426_o;
  wire n5428_o;
  wire n5430_o;
  wire n5432_o;
  wire n5433_o;
  wire n5435_o;
  wire n5437_o;
  wire [1:0] n5438_o;
  wire [3:0] n5439_o;
  wire [1:0] n5440_o;
  wire n5441_o;
  wire n5442_o;
  wire n5443_o;
  wire n5444_o;
  wire n5445_o;
  wire n5446_o;
  wire n5447_o;
  wire n5448_o;
  wire n5449_o;
  wire n5450_o;
  wire n5451_o;
  wire n5452_o;
  wire n5453_o;
  wire n5454_o;
  wire n5455_o;
  wire n5456_o;
  wire n5457_o;
  wire n5458_o;
  wire n5459_o;
  wire [3:0] n5460_o;
  wire [3:0] n5461_o;
  wire n5462_o;
  wire [1:0] n5463_o;
  wire n5464_o;
  wire n5465_o;
  wire [2:0] n5466_o;
  wire n5468_o;
  wire n5470_o;
  wire [2:0] n5472_o;
  wire [6:0] n5473_o;
  wire n5475_o;
  wire [6:0] n5476_o;
  reg n5477_o;
  reg [1:0] n5478_o;
  reg [1:0] n5479_o;
  reg n5480_o;
  reg n5481_o;
  reg n5483_o;
  reg n5484_o;
  reg n5486_o;
  reg n5488_o;
  reg n5490_o;
  reg n5492_o;
  reg n5494_o;
  reg n5496_o;
  reg n5498_o;
  reg n5500_o;
  reg [5:0] n5501_o;
  reg n5503_o;
  reg n5504_o;
  reg n5506_o;
  reg n5508_o;
  reg n5510_o;
  reg n5512_o;
  reg n5514_o;
  reg n5516_o;
  reg n5518_o;
  wire n5519_o;
  reg n5520_o;
  wire n5521_o;
  reg n5522_o;
  wire n5523_o;
  reg n5524_o;
  wire n5525_o;
  reg n5526_o;
  wire n5527_o;
  reg n5528_o;
  wire n5529_o;
  reg n5530_o;
  wire n5531_o;
  reg n5532_o;
  wire n5533_o;
  wire n5534_o;
  wire n5535_o;
  reg n5536_o;
  wire n5537_o;
  wire n5538_o;
  wire n5539_o;
  reg n5540_o;
  wire n5541_o;
  reg n5542_o;
  wire n5543_o;
  reg n5544_o;
  wire n5545_o;
  wire n5546_o;
  reg n5547_o;
  wire n5548_o;
  wire n5549_o;
  reg n5550_o;
  wire n5551_o;
  reg n5552_o;
  wire n5553_o;
  reg n5554_o;
  wire n5555_o;
  reg n5556_o;
  wire n5557_o;
  reg n5558_o;
  wire [3:0] n5559_o;
  reg [3:0] n5560_o;
  reg [1:0] n5561_o;
  reg [1:0] n5562_o;
  wire n5563_o;
  reg n5564_o;
  wire n5565_o;
  reg n5566_o;
  reg n5567_o;
  wire n5568_o;
  reg n5569_o;
  reg n5571_o;
  wire n5572_o;
  reg n5574_o;
  wire n5575_o;
  reg n5577_o;
  reg n5579_o;
  reg n5581_o;
  reg n5583_o;
  reg n5585_o;
  reg n5587_o;
  reg n5589_o;
  reg n5591_o;
  reg n5593_o;
  wire [1:0] n5594_o;
  reg [1:0] n5596_o;
  wire n5597_o;
  reg n5599_o;
  reg n5601_o;
  reg [6:0] n5602_o;
  wire n5603_o;
  wire [1:0] n5604_o;
  wire [1:0] n5605_o;
  wire n5606_o;
  wire n5607_o;
  wire n5609_o;
  wire n5610_o;
  wire n5612_o;
  wire n5614_o;
  wire n5615_o;
  wire n5616_o;
  wire n5617_o;
  wire n5619_o;
  wire n5621_o;
  wire n5623_o;
  wire n5624_o;
  wire [5:0] n5625_o;
  wire n5627_o;
  wire n5628_o;
  wire n5629_o;
  wire n5631_o;
  wire n5633_o;
  wire n5635_o;
  wire n5636_o;
  wire n5638_o;
  wire n5639_o;
  wire [3:0] n5640_o;
  wire [9:0] n5641_o;
  wire [3:0] n5642_o;
  wire [1:0] n5643_o;
  wire n5644_o;
  wire n5645_o;
  wire n5646_o;
  wire n5647_o;
  wire n5648_o;
  wire n5649_o;
  wire n5650_o;
  wire n5651_o;
  wire n5652_o;
  wire n5653_o;
  wire n5654_o;
  wire n5655_o;
  wire n5656_o;
  wire n5657_o;
  wire n5658_o;
  wire n5659_o;
  wire [2:0] n5660_o;
  wire n5661_o;
  wire [2:0] n5662_o;
  wire [2:0] n5663_o;
  wire n5664_o;
  wire n5665_o;
  wire [4:0] n5666_o;
  wire [4:0] n5667_o;
  wire [4:0] n5668_o;
  wire n5669_o;
  wire n5670_o;
  wire [3:0] n5671_o;
  wire [3:0] n5672_o;
  wire [3:0] n5673_o;
  wire [3:0] n5674_o;
  wire [3:0] n5675_o;
  wire n5676_o;
  wire n5677_o;
  wire n5678_o;
  wire n5679_o;
  wire n5680_o;
  wire [1:0] n5681_o;
  wire [1:0] n5682_o;
  wire [1:0] n5683_o;
  wire [1:0] n5684_o;
  wire [2:0] n5685_o;
  wire n5686_o;
  wire [1:0] n5688_o;
  wire [1:0] n5690_o;
  wire n5691_o;
  wire n5693_o;
  wire n5695_o;
  wire n5697_o;
  wire n5699_o;
  wire n5701_o;
  wire n5703_o;
  wire [1:0] n5704_o;
  wire [1:0] n5706_o;
  wire n5707_o;
  wire n5708_o;
  wire n5709_o;
  wire [6:0] n5710_o;
  wire n5712_o;
  wire [1:0] n5713_o;
  wire n5715_o;
  wire [2:0] n5716_o;
  wire n5718_o;
  wire n5722_o;
  wire n5723_o;
  wire n5724_o;
  wire [6:0] n5726_o;
  wire [2:0] n5727_o;
  wire n5729_o;
  wire [1:0] n5730_o;
  wire n5732_o;
  wire [2:0] n5733_o;
  wire n5735_o;
  wire n5736_o;
  wire n5737_o;
  wire n5738_o;
  wire [1:0] n5739_o;
  wire n5741_o;
  wire n5742_o;
  wire n5744_o;
  wire n5745_o;
  wire [6:0] n5747_o;
  wire [1:0] n5749_o;
  wire [1:0] n5750_o;
  wire n5751_o;
  wire n5752_o;
  wire n5753_o;
  wire n5754_o;
  wire n5757_o;
  wire n5760_o;
  wire [1:0] n5761_o;
  wire n5764_o;
  wire n5766_o;
  wire n5768_o;
  wire n5769_o;
  wire n5770_o;
  wire [2:0] n5771_o;
  wire n5773_o;
  wire [1:0] n5774_o;
  wire n5776_o;
  wire n5777_o;
  wire n5779_o;
  wire n5781_o;
  wire n5782_o;
  wire n5783_o;
  wire n5784_o;
  wire n5786_o;
  wire [1:0] n5787_o;
  wire n5789_o;
  wire n5792_o;
  wire n5793_o;
  wire [1:0] n5795_o;
  wire n5798_o;
  wire n5801_o;
  wire n5804_o;
  wire n5807_o;
  wire n5809_o;
  wire n5811_o;
  wire n5812_o;
  wire [1:0] n5813_o;
  wire n5814_o;
  wire n5816_o;
  wire n5817_o;
  wire n5819_o;
  wire n5820_o;
  wire n5822_o;
  wire n5823_o;
  wire n5825_o;
  wire n5827_o;
  wire n5828_o;
  wire n5829_o;
  wire [1:0] n5830_o;
  wire [1:0] n5831_o;
  wire n5833_o;
  wire n5835_o;
  wire n5837_o;
  wire n5839_o;
  wire n5841_o;
  wire n5843_o;
  wire n5845_o;
  wire n5846_o;
  wire n5848_o;
  wire n5850_o;
  wire [6:0] n5851_o;
  wire [4:0] n5852_o;
  wire n5854_o;
  wire [2:0] n5855_o;
  wire n5857_o;
  wire [1:0] n5858_o;
  wire n5860_o;
  wire n5861_o;
  wire n5862_o;
  wire [2:0] n5863_o;
  wire n5865_o;
  wire n5867_o;
  wire n5868_o;
  wire n5869_o;
  wire n5871_o;
  wire n5872_o;
  wire [1:0] n5876_o;
  wire n5878_o;
  wire n5881_o;
  wire n5884_o;
  wire n5887_o;
  wire n5890_o;
  wire n5893_o;
  wire n5895_o;
  wire n5897_o;
  wire [1:0] n5898_o;
  wire [1:0] n5900_o;
  wire n5902_o;
  wire n5904_o;
  wire n5905_o;
  wire [1:0] n5906_o;
  wire [1:0] n5907_o;
  wire n5909_o;
  wire n5910_o;
  wire n5911_o;
  wire n5913_o;
  wire n5914_o;
  wire n5915_o;
  wire n5916_o;
  wire n5917_o;
  wire n5919_o;
  wire n5920_o;
  wire n5921_o;
  wire n5922_o;
  wire [1:0] n5924_o;
  wire n5926_o;
  wire n5928_o;
  wire n5929_o;
  wire [6:0] n5930_o;
  wire n5932_o;
  wire n5934_o;
  wire [3:0] n5935_o;
  wire n5937_o;
  wire [7:0] n5939_o;
  wire n5941_o;
  wire [7:0] n5943_o;
  wire n5945_o;
  wire [1:0] n5947_o;
  wire n5950_o;
  wire [6:0] n5953_o;
  wire [1:0] n5954_o;
  wire n5956_o;
  wire n5957_o;
  wire [6:0] n5959_o;
  wire [7:0] n5960_o;
  wire n5962_o;
  wire [7:0] n5964_o;
  wire n5966_o;
  wire [1:0] n5968_o;
  wire [1:0] n5969_o;
  wire n5970_o;
  wire [1:0] n5971_o;
  wire n5973_o;
  wire n5975_o;
  wire n5976_o;
  wire n5977_o;
  wire n5978_o;
  wire n5979_o;
  wire n5980_o;
  wire [6:0] n5982_o;
  wire [1:0] n5983_o;
  wire n5984_o;
  wire n5986_o;
  wire n5987_o;
  wire n5988_o;
  wire n5989_o;
  wire n5990_o;
  wire n5991_o;
  wire [6:0] n5992_o;
  wire n5994_o;
  wire n5995_o;
  wire n5996_o;
  wire [1:0] n6001_o;
  wire n6004_o;
  wire n6007_o;
  wire n6010_o;
  wire [1:0] n6011_o;
  wire [1:0] n6013_o;
  wire n6015_o;
  wire n6017_o;
  wire [1:0] n6018_o;
  wire n6020_o;
  wire [2:0] n6021_o;
  wire n6023_o;
  wire n6025_o;
  wire [3:0] n6026_o;
  wire n6028_o;
  wire [1:0] n6029_o;
  wire n6031_o;
  wire n6032_o;
  wire n6033_o;
  wire [1:0] n6034_o;
  wire n6036_o;
  wire n6039_o;
  wire n6041_o;
  wire n6042_o;
  wire [1:0] n6043_o;
  wire n6045_o;
  wire n6046_o;
  wire n6047_o;
  wire [1:0] n6049_o;
  wire [6:0] n6051_o;
  wire n6052_o;
  wire n6053_o;
  wire n6054_o;
  wire n6057_o;
  wire [1:0] n6058_o;
  wire n6060_o;
  wire n6061_o;
  wire n6062_o;
  wire n6065_o;
  wire [1:0] n6067_o;
  wire n6068_o;
  wire n6070_o;
  wire n6073_o;
  wire n6075_o;
  wire n6078_o;
  wire n6081_o;
  wire n6084_o;
  wire n6086_o;
  wire n6087_o;
  wire n6088_o;
  wire [1:0] n6089_o;
  wire n6091_o;
  wire n6092_o;
  wire [1:0] n6093_o;
  wire n6095_o;
  wire [1:0] n6099_o;
  wire n6101_o;
  wire [1:0] n6102_o;
  wire n6104_o;
  wire n6105_o;
  wire [1:0] n6108_o;
  wire n6110_o;
  wire [1:0] n6115_o;
  wire n6117_o;
  wire n6119_o;
  wire n6120_o;
  wire n6121_o;
  wire [1:0] n6122_o;
  wire n6124_o;
  wire [1:0] n6127_o;
  wire n6131_o;
  wire n6132_o;
  wire n6133_o;
  wire n6134_o;
  wire [6:0] n6136_o;
  wire n6138_o;
  wire [6:0] n6140_o;
  wire [1:0] n6141_o;
  wire n6144_o;
  wire n6147_o;
  wire n6148_o;
  wire n6150_o;
  wire n6152_o;
  wire n6154_o;
  wire [6:0] n6155_o;
  wire [1:0] n6156_o;
  wire n6157_o;
  wire n6159_o;
  wire n6162_o;
  wire n6164_o;
  wire n6165_o;
  wire n6168_o;
  wire n6171_o;
  wire n6173_o;
  wire n6174_o;
  wire n6175_o;
  wire n6177_o;
  wire [1:0] n6178_o;
  wire n6180_o;
  wire n6182_o;
  wire [1:0] n6184_o;
  wire [6:0] n6185_o;
  wire [1:0] n6186_o;
  wire [1:0] n6187_o;
  wire n6189_o;
  wire n6191_o;
  wire n6193_o;
  wire n6194_o;
  wire n6196_o;
  wire n6198_o;
  wire n6201_o;
  wire n6202_o;
  wire n6203_o;
  wire n6204_o;
  wire n6205_o;
  wire n6206_o;
  wire n6207_o;
  wire n6208_o;
  wire n6209_o;
  wire n6211_o;
  wire n6213_o;
  wire n6215_o;
  wire n6217_o;
  wire [1:0] n6219_o;
  wire [6:0] n6220_o;
  wire [1:0] n6221_o;
  wire n6223_o;
  wire n6224_o;
  wire n6225_o;
  wire [2:0] n6226_o;
  wire n6228_o;
  wire n6229_o;
  wire [3:0] n6230_o;
  wire n6232_o;
  wire [1:0] n6233_o;
  wire n6235_o;
  wire n6236_o;
  wire n6237_o;
  wire n6238_o;
  wire [1:0] n6239_o;
  wire n6241_o;
  wire n6242_o;
  wire [2:0] n6243_o;
  wire n6245_o;
  wire [1:0] n6246_o;
  wire n6248_o;
  wire n6249_o;
  wire n6250_o;
  wire n6251_o;
  wire n6252_o;
  wire n6256_o;
  wire n6259_o;
  wire n6262_o;
  wire n6264_o;
  wire [1:0] n6265_o;
  wire [1:0] n6266_o;
  wire n6268_o;
  wire n6270_o;
  wire n6272_o;
  wire n6273_o;
  wire n6274_o;
  wire n6275_o;
  wire n6277_o;
  wire n6279_o;
  wire n6280_o;
  wire n6281_o;
  wire n6282_o;
  wire n6283_o;
  wire n6285_o;
  wire n6286_o;
  wire n6287_o;
  wire n6289_o;
  wire n6291_o;
  wire n6293_o;
  wire n6295_o;
  wire n6297_o;
  wire [1:0] n6299_o;
  wire [6:0] n6300_o;
  wire [1:0] n6301_o;
  wire [1:0] n6302_o;
  wire n6303_o;
  wire n6305_o;
  wire n6307_o;
  wire n6308_o;
  wire n6309_o;
  wire n6310_o;
  wire n6311_o;
  wire n6312_o;
  wire n6314_o;
  wire n6316_o;
  wire n6318_o;
  wire n6319_o;
  wire n6320_o;
  wire n6321_o;
  wire n6322_o;
  wire n6323_o;
  wire n6324_o;
  wire n6325_o;
  wire n6326_o;
  wire n6328_o;
  wire n6330_o;
  wire n6332_o;
  wire n6334_o;
  wire n6335_o;
  wire [1:0] n6337_o;
  wire [6:0] n6338_o;
  wire n6340_o;
  wire [5:0] n6341_o;
  wire n6343_o;
  wire n6344_o;
  wire n6345_o;
  wire [1:0] n6346_o;
  wire n6348_o;
  wire n6349_o;
  wire [3:0] n6350_o;
  wire n6352_o;
  wire [1:0] n6353_o;
  wire n6355_o;
  wire n6356_o;
  wire n6357_o;
  wire n6358_o;
  wire [2:0] n6359_o;
  wire n6361_o;
  wire [1:0] n6362_o;
  wire n6364_o;
  wire n6365_o;
  wire n6366_o;
  wire n6367_o;
  wire n6368_o;
  wire n6370_o;
  wire n6371_o;
  wire n6373_o;
  wire n6374_o;
  wire [1:0] n6375_o;
  wire n6377_o;
  wire n6378_o;
  wire n6379_o;
  wire [1:0] n6381_o;
  wire n6383_o;
  wire n6386_o;
  wire n6390_o;
  wire n6393_o;
  wire n6394_o;
  wire [1:0] n6395_o;
  wire n6397_o;
  wire n6398_o;
  wire n6401_o;
  wire n6404_o;
  wire n6405_o;
  wire n6407_o;
  wire n6410_o;
  wire n6412_o;
  wire n6414_o;
  wire n6416_o;
  wire n6418_o;
  wire n6419_o;
  wire n6420_o;
  wire n6422_o;
  wire n6423_o;
  wire n6425_o;
  wire n6427_o;
  wire n6429_o;
  wire n6431_o;
  wire n6434_o;
  wire n6437_o;
  wire n6440_o;
  wire n6442_o;
  wire n6444_o;
  wire n6446_o;
  wire n6448_o;
  wire n6450_o;
  wire n6452_o;
  wire n6454_o;
  wire n6456_o;
  wire n6457_o;
  wire n6459_o;
  wire [1:0] n6460_o;
  wire n6462_o;
  wire [3:0] n6463_o;
  wire n6465_o;
  wire [1:0] n6466_o;
  wire n6468_o;
  wire n6469_o;
  wire n6470_o;
  wire n6471_o;
  wire [1:0] n6474_o;
  wire n6476_o;
  wire n6478_o;
  wire n6481_o;
  wire n6483_o;
  wire n6486_o;
  wire n6489_o;
  wire n6492_o;
  wire n6494_o;
  wire n6496_o;
  wire n6498_o;
  wire n6500_o;
  wire n6502_o;
  wire n6505_o;
  wire n6508_o;
  wire n6511_o;
  wire n6512_o;
  wire n6513_o;
  wire n6515_o;
  wire n6517_o;
  wire n6518_o;
  wire [2:0] n6519_o;
  wire n6521_o;
  wire [2:0] n6523_o;
  wire n6525_o;
  wire n6527_o;
  wire [1:0] n6531_o;
  wire n6532_o;
  wire n6533_o;
  wire n6534_o;
  wire n6535_o;
  wire n6536_o;
  wire n6537_o;
  wire [6:0] n6539_o;
  wire [2:0] n6542_o;
  wire n6544_o;
  wire [1:0] n6545_o;
  wire n6547_o;
  wire n6548_o;
  wire n6552_o;
  wire n6555_o;
  wire n6558_o;
  wire n6561_o;
  wire n6563_o;
  wire n6564_o;
  wire n6566_o;
  wire n6568_o;
  wire n6570_o;
  wire n6572_o;
  wire n6573_o;
  wire n6574_o;
  wire n6575_o;
  wire n6576_o;
  wire n6577_o;
  wire n6578_o;
  wire n6579_o;
  wire n6580_o;
  wire n6582_o;
  wire n6584_o;
  wire n6586_o;
  wire n6587_o;
  wire [5:0] n6588_o;
  wire n6590_o;
  wire [3:0] n6591_o;
  wire n6593_o;
  wire [1:0] n6594_o;
  wire n6596_o;
  wire n6597_o;
  wire n6598_o;
  wire n6603_o;
  wire n6606_o;
  wire n6609_o;
  wire n6612_o;
  wire n6613_o;
  wire n6614_o;
  wire n6616_o;
  wire n6617_o;
  wire n6618_o;
  wire n6619_o;
  wire n6620_o;
  wire n6621_o;
  wire n6622_o;
  wire n6623_o;
  wire n6624_o;
  wire n6625_o;
  wire n6626_o;
  wire n6627_o;
  wire n6628_o;
  wire [1:0] n6629_o;
  wire n6630_o;
  wire n6632_o;
  wire n6633_o;
  wire n6634_o;
  wire n6636_o;
  wire n6637_o;
  wire n6638_o;
  wire [1:0] n6639_o;
  wire n6641_o;
  wire n6643_o;
  wire n6645_o;
  wire n6647_o;
  wire n6648_o;
  wire n6649_o;
  wire n6650_o;
  wire n6652_o;
  wire n6653_o;
  wire n6654_o;
  wire n6655_o;
  wire n6656_o;
  wire n6657_o;
  wire n6658_o;
  wire n6659_o;
  wire [1:0] n6660_o;
  wire n6661_o;
  wire n6663_o;
  wire n6664_o;
  wire n6665_o;
  wire n6667_o;
  wire n6669_o;
  wire [6:0] n6670_o;
  wire n6672_o;
  wire [1:0] n6673_o;
  wire n6675_o;
  wire [2:0] n6676_o;
  wire n6678_o;
  wire n6680_o;
  wire [3:0] n6681_o;
  wire n6683_o;
  wire [1:0] n6684_o;
  wire n6686_o;
  wire n6687_o;
  wire n6688_o;
  wire [1:0] n6689_o;
  wire n6691_o;
  wire n6694_o;
  wire n6696_o;
  wire n6697_o;
  wire [1:0] n6698_o;
  wire n6700_o;
  wire n6701_o;
  wire n6702_o;
  wire [1:0] n6705_o;
  wire n6706_o;
  wire n6707_o;
  wire [6:0] n6709_o;
  wire [1:0] n6711_o;
  wire n6713_o;
  wire n6714_o;
  wire n6715_o;
  wire n6718_o;
  wire [1:0] n6721_o;
  wire [1:0] n6723_o;
  wire n6724_o;
  wire n6726_o;
  wire n6729_o;
  wire n6731_o;
  wire n6734_o;
  wire n6737_o;
  wire n6740_o;
  wire n6742_o;
  wire n6744_o;
  wire n6745_o;
  wire n6746_o;
  wire [1:0] n6747_o;
  wire n6749_o;
  wire n6750_o;
  wire [1:0] n6751_o;
  wire n6753_o;
  wire [3:0] n6756_o;
  wire n6758_o;
  wire [4:0] n6759_o;
  wire n6761_o;
  wire n6762_o;
  wire n6766_o;
  wire n6767_o;
  wire n6768_o;
  wire n6771_o;
  wire n6774_o;
  wire [1:0] n6776_o;
  wire n6779_o;
  wire [1:0] n6781_o;
  wire n6782_o;
  wire n6784_o;
  wire n6786_o;
  wire n6788_o;
  wire n6791_o;
  wire n6794_o;
  wire n6795_o;
  wire n6796_o;
  wire n6797_o;
  wire n6798_o;
  wire n6799_o;
  wire n6800_o;
  wire [1:0] n6801_o;
  wire [1:0] n6802_o;
  wire n6804_o;
  wire n6806_o;
  wire n6808_o;
  wire n6810_o;
  wire n6812_o;
  wire n6815_o;
  wire n6816_o;
  wire n6817_o;
  wire n6818_o;
  wire n6819_o;
  wire n6820_o;
  wire n6821_o;
  wire n6823_o;
  wire n6825_o;
  wire [1:0] n6826_o;
  wire n6828_o;
  wire n6829_o;
  wire n6830_o;
  wire [2:0] n6831_o;
  wire n6833_o;
  wire n6834_o;
  wire [3:0] n6835_o;
  wire n6837_o;
  wire [1:0] n6838_o;
  wire n6840_o;
  wire n6841_o;
  wire n6842_o;
  wire n6843_o;
  wire [1:0] n6844_o;
  wire n6846_o;
  wire n6847_o;
  wire [2:0] n6848_o;
  wire n6850_o;
  wire [1:0] n6851_o;
  wire n6853_o;
  wire n6854_o;
  wire n6855_o;
  wire n6856_o;
  wire n6857_o;
  wire n6861_o;
  wire n6864_o;
  wire n6867_o;
  wire n6869_o;
  wire [1:0] n6870_o;
  wire [1:0] n6871_o;
  wire n6873_o;
  wire n6875_o;
  wire n6877_o;
  wire n6878_o;
  wire n6879_o;
  wire n6881_o;
  wire n6883_o;
  wire n6884_o;
  wire n6885_o;
  wire n6886_o;
  wire n6887_o;
  wire n6888_o;
  wire n6889_o;
  wire n6891_o;
  wire n6893_o;
  wire n6895_o;
  wire [1:0] n6896_o;
  wire [1:0] n6897_o;
  wire n6899_o;
  wire n6901_o;
  wire n6903_o;
  wire n6905_o;
  wire n6906_o;
  wire n6907_o;
  wire n6908_o;
  wire n6910_o;
  wire n6912_o;
  wire n6914_o;
  wire n6916_o;
  wire n6917_o;
  wire n6918_o;
  wire n6919_o;
  wire n6920_o;
  wire n6921_o;
  wire n6922_o;
  wire n6924_o;
  wire n6926_o;
  wire n6928_o;
  wire n6930_o;
  wire n6931_o;
  wire n6933_o;
  wire [1:0] n6934_o;
  wire n6936_o;
  wire n6937_o;
  wire n6938_o;
  wire [1:0] n6939_o;
  wire n6941_o;
  wire [2:0] n6942_o;
  wire n6944_o;
  wire [1:0] n6945_o;
  wire n6947_o;
  wire n6948_o;
  wire n6949_o;
  wire [1:0] n6951_o;
  wire [1:0] n6954_o;
  wire n6957_o;
  wire [1:0] n6958_o;
  wire n6961_o;
  wire n6964_o;
  wire n6967_o;
  wire n6969_o;
  wire n6971_o;
  wire n6972_o;
  wire n6973_o;
  wire n6975_o;
  wire n6977_o;
  wire [1:0] n6978_o;
  wire n6980_o;
  wire [2:0] n6981_o;
  wire n6983_o;
  wire n6984_o;
  wire [2:0] n6985_o;
  wire n6987_o;
  wire n6988_o;
  wire [2:0] n6989_o;
  wire n6991_o;
  wire [2:0] n6992_o;
  wire n6994_o;
  wire n6995_o;
  wire [2:0] n6996_o;
  wire n6998_o;
  wire n6999_o;
  wire [2:0] n7000_o;
  wire n7002_o;
  wire [1:0] n7003_o;
  wire n7005_o;
  wire n7006_o;
  wire n7007_o;
  wire n7008_o;
  wire n7009_o;
  wire [1:0] n7010_o;
  wire n7012_o;
  wire [2:0] n7013_o;
  wire n7015_o;
  wire n7016_o;
  wire [2:0] n7017_o;
  wire n7019_o;
  wire n7020_o;
  wire [2:0] n7021_o;
  wire n7023_o;
  wire [2:0] n7024_o;
  wire n7026_o;
  wire n7027_o;
  wire [2:0] n7028_o;
  wire n7030_o;
  wire n7031_o;
  wire [3:0] n7032_o;
  wire n7034_o;
  wire n7035_o;
  wire n7036_o;
  wire n7037_o;
  wire n7040_o;
  wire n7041_o;
  wire n7042_o;
  wire n7043_o;
  wire [6:0] n7045_o;
  wire n7047_o;
  wire n7048_o;
  wire n7049_o;
  wire n7050_o;
  wire n7053_o;
  wire [2:0] n7054_o;
  wire n7056_o;
  wire n7059_o;
  wire [2:0] n7060_o;
  wire n7062_o;
  wire [2:0] n7063_o;
  wire n7065_o;
  wire n7066_o;
  wire [2:0] n7067_o;
  wire n7069_o;
  wire n7070_o;
  wire [2:0] n7071_o;
  wire n7073_o;
  wire n7074_o;
  wire n7077_o;
  wire [2:0] n7078_o;
  wire n7080_o;
  wire [2:0] n7081_o;
  wire n7083_o;
  wire n7084_o;
  wire [2:0] n7085_o;
  wire n7087_o;
  wire n7088_o;
  wire n7091_o;
  wire [1:0] n7092_o;
  wire n7094_o;
  wire [2:0] n7095_o;
  wire n7097_o;
  wire n7099_o;
  wire n7100_o;
  wire [1:0] n7103_o;
  wire n7106_o;
  wire n7109_o;
  wire n7110_o;
  wire n7111_o;
  wire n7112_o;
  wire n7114_o;
  wire n7116_o;
  wire n7118_o;
  wire n7119_o;
  wire n7120_o;
  wire [1:0] n7122_o;
  wire n7123_o;
  wire [1:0] n7127_o;
  wire n7129_o;
  wire n7131_o;
  wire n7132_o;
  wire n7133_o;
  wire n7134_o;
  wire [6:0] n7136_o;
  wire [2:0] n7137_o;
  wire n7139_o;
  wire n7142_o;
  wire n7145_o;
  wire [2:0] n7146_o;
  wire n7148_o;
  wire [2:0] n7149_o;
  wire n7151_o;
  wire n7152_o;
  wire [2:0] n7153_o;
  wire n7155_o;
  wire n7156_o;
  wire n7158_o;
  wire n7160_o;
  wire n7162_o;
  wire n7163_o;
  wire [1:0] n7164_o;
  wire n7166_o;
  wire n7169_o;
  wire n7171_o;
  wire n7173_o;
  wire n7175_o;
  wire n7177_o;
  wire n7180_o;
  wire n7183_o;
  wire n7184_o;
  wire n7185_o;
  wire n7186_o;
  wire n7187_o;
  wire n7188_o;
  wire n7189_o;
  wire n7190_o;
  wire n7191_o;
  wire [1:0] n7192_o;
  wire n7194_o;
  wire n7196_o;
  wire [1:0] n7198_o;
  wire [6:0] n7199_o;
  wire n7200_o;
  wire [1:0] n7201_o;
  wire n7202_o;
  wire n7204_o;
  wire n7206_o;
  wire n7208_o;
  wire n7210_o;
  wire n7212_o;
  wire n7213_o;
  wire n7214_o;
  wire n7215_o;
  wire n7217_o;
  wire n7218_o;
  wire n7219_o;
  wire n7220_o;
  wire n7221_o;
  wire n7222_o;
  wire n7223_o;
  wire n7224_o;
  wire n7225_o;
  wire n7227_o;
  wire n7228_o;
  wire n7230_o;
  wire [1:0] n7232_o;
  wire [6:0] n7233_o;
  wire n7237_o;
  wire [2:0] n7239_o;
  wire [2:0] n7240_o;
  wire n7242_o;
  wire n7245_o;
  wire [1:0] n7247_o;
  wire [3:0] n7248_o;
  wire [3:0] n7249_o;
  wire [3:0] n7250_o;
  wire [3:0] n7251_o;
  wire [3:0] n7252_o;
  wire n7253_o;
  wire n7254_o;
  wire [6:0] n7256_o;
  wire n7257_o;
  wire [3:0] n7258_o;
  wire [3:0] n7259_o;
  wire [3:0] n7260_o;
  wire [3:0] n7261_o;
  wire n7263_o;
  wire n7264_o;
  wire n7265_o;
  wire [1:0] n7266_o;
  wire n7269_o;
  wire n7271_o;
  wire n7273_o;
  wire n7275_o;
  wire n7277_o;
  wire n7279_o;
  wire n7281_o;
  wire n7282_o;
  wire [3:0] n7283_o;
  wire [3:0] n7284_o;
  wire [3:0] n7285_o;
  wire [3:0] n7286_o;
  wire n7288_o;
  wire n7290_o;
  wire n7292_o;
  wire n7293_o;
  wire n7294_o;
  wire n7295_o;
  wire n7296_o;
  wire n7297_o;
  wire n7298_o;
  wire n7299_o;
  wire n7300_o;
  wire n7301_o;
  wire n7302_o;
  wire n7303_o;
  wire n7305_o;
  wire n7306_o;
  wire [1:0] n7308_o;
  wire [6:0] n7309_o;
  wire n7311_o;
  wire n7312_o;
  wire [2:0] n7313_o;
  wire n7315_o;
  wire n7316_o;
  wire [1:0] n7317_o;
  wire n7319_o;
  wire [2:0] n7320_o;
  wire n7322_o;
  wire n7323_o;
  wire [2:0] n7324_o;
  wire n7326_o;
  wire [1:0] n7327_o;
  wire n7329_o;
  wire n7330_o;
  wire n7331_o;
  wire [2:0] n7332_o;
  wire n7334_o;
  wire n7335_o;
  wire n7336_o;
  wire [1:0] n7337_o;
  wire n7339_o;
  wire n7340_o;
  wire n7343_o;
  wire n7346_o;
  wire n7348_o;
  wire n7351_o;
  wire n7353_o;
  wire n7356_o;
  wire n7359_o;
  wire n7361_o;
  wire n7362_o;
  wire n7363_o;
  wire n7365_o;
  wire n7367_o;
  wire n7369_o;
  wire n7370_o;
  wire [2:0] n7371_o;
  wire n7373_o;
  wire n7374_o;
  wire [1:0] n7375_o;
  wire n7377_o;
  wire [2:0] n7378_o;
  wire n7380_o;
  wire n7381_o;
  wire [2:0] n7382_o;
  wire n7384_o;
  wire [1:0] n7385_o;
  wire n7387_o;
  wire [2:0] n7388_o;
  wire n7390_o;
  wire n7391_o;
  wire n7392_o;
  wire n7393_o;
  wire [4:0] n7394_o;
  wire n7396_o;
  wire [2:0] n7397_o;
  wire n7399_o;
  wire [2:0] n7400_o;
  wire n7402_o;
  wire n7403_o;
  wire [2:0] n7404_o;
  wire n7406_o;
  wire n7409_o;
  wire n7412_o;
  wire n7414_o;
  wire n7417_o;
  wire n7419_o;
  wire n7422_o;
  wire n7425_o;
  wire n7427_o;
  wire n7428_o;
  wire n7429_o;
  wire n7431_o;
  wire n7433_o;
  wire n7435_o;
  wire n7437_o;
  wire n7439_o;
  wire n7441_o;
  wire n7443_o;
  wire n7445_o;
  wire n7447_o;
  wire n7448_o;
  wire n7449_o;
  wire n7450_o;
  wire n7452_o;
  wire [12:0] n7453_o;
  reg n7454_o;
  reg [1:0] n7456_o;
  reg [1:0] n7457_o;
  reg [1:0] n7458_o;
  reg n7459_o;
  reg n7461_o;
  reg n7462_o;
  reg n7464_o;
  reg n7466_o;
  reg n7467_o;
  reg n7469_o;
  reg n7471_o;
  reg n7473_o;
  reg n7475_o;
  reg n7477_o;
  reg n7479_o;
  reg n7481_o;
  reg n7483_o;
  reg n7485_o;
  reg n7487_o;
  reg [1:0] n7488_o;
  wire [3:0] n7489_o;
  wire [3:0] n7490_o;
  wire [3:0] n7491_o;
  wire [3:0] n7492_o;
  reg [3:0] n7493_o;
  wire [1:0] n7494_o;
  wire [1:0] n7495_o;
  wire [1:0] n7496_o;
  wire [1:0] n7497_o;
  reg [1:0] n7498_o;
  reg n7500_o;
  reg n7501_o;
  reg n7504_o;
  reg n7506_o;
  reg n7509_o;
  reg n7511_o;
  reg n7513_o;
  reg n7515_o;
  reg n7520_o;
  reg n7522_o;
  reg n7524_o;
  reg n7526_o;
  reg n7528_o;
  reg n7530_o;
  wire n7531_o;
  reg n7532_o;
  wire [2:0] n7533_o;
  reg [2:0] n7534_o;
  wire n7535_o;
  reg n7536_o;
  wire n7537_o;
  reg n7538_o;
  wire n7539_o;
  reg n7540_o;
  wire n7541_o;
  reg n7542_o;
  wire n7543_o;
  reg n7544_o;
  wire n7545_o;
  reg n7546_o;
  reg n7547_o;
  wire n7548_o;
  reg n7549_o;
  wire n7550_o;
  reg n7551_o;
  wire n7552_o;
  wire n7553_o;
  reg n7554_o;
  wire n7555_o;
  wire n7556_o;
  reg n7557_o;
  wire n7558_o;
  reg n7559_o;
  wire n7560_o;
  wire n7561_o;
  wire n7562_o;
  wire n7563_o;
  wire n7564_o;
  reg n7565_o;
  wire n7566_o;
  wire n7567_o;
  wire n7568_o;
  wire n7569_o;
  wire n7570_o;
  reg n7571_o;
  wire n7572_o;
  wire n7573_o;
  reg n7574_o;
  wire n7575_o;
  wire n7576_o;
  reg n7577_o;
  wire n7578_o;
  reg n7579_o;
  wire [1:0] n7580_o;
  wire [1:0] n7581_o;
  reg [1:0] n7582_o;
  wire n7583_o;
  wire n7584_o;
  reg n7585_o;
  wire n7586_o;
  wire n7587_o;
  reg n7588_o;
  wire n7589_o;
  wire n7590_o;
  wire n7591_o;
  reg n7592_o;
  wire n7593_o;
  wire n7594_o;
  reg n7595_o;
  wire [3:0] n7596_o;
  reg [3:0] n7597_o;
  wire n7598_o;
  reg n7599_o;
  wire [3:0] n7600_o;
  reg [3:0] n7601_o;
  wire n7602_o;
  reg n7603_o;
  wire n7604_o;
  reg n7605_o;
  wire n7606_o;
  reg n7607_o;
  wire n7608_o;
  wire n7609_o;
  reg n7610_o;
  wire n7611_o;
  reg n7612_o;
  wire n7613_o;
  reg n7614_o;
  wire n7615_o;
  reg n7616_o;
  wire n7617_o;
  reg n7618_o;
  wire n7619_o;
  reg n7620_o;
  wire n7621_o;
  reg n7623_o;
  wire n7624_o;
  reg n7626_o;
  wire n7627_o;
  reg n7629_o;
  wire n7630_o;
  wire n7631_o;
  reg n7633_o;
  wire n7634_o;
  reg n7636_o;
  wire n7637_o;
  reg n7639_o;
  wire n7640_o;
  wire n7641_o;
  reg n7643_o;
  wire n7644_o;
  wire n7645_o;
  reg n7647_o;
  wire n7648_o;
  reg n7650_o;
  reg n7652_o;
  reg n7654_o;
  reg n7656_o;
  reg n7658_o;
  reg n7660_o;
  reg n7662_o;
  reg n7664_o;
  reg n7666_o;
  reg n7668_o;
  reg n7670_o;
  reg n7672_o;
  reg n7674_o;
  reg [1:0] n7676_o;
  reg n7678_o;
  reg [1:0] n7680_o;
  reg [1:0] n7682_o;
  reg n7684_o;
  reg [6:0] n7685_o;
  wire n7686_o;
  wire [1:0] n7687_o;
  wire [1:0] n7688_o;
  wire [1:0] n7689_o;
  wire n7690_o;
  wire n7692_o;
  wire n7694_o;
  wire n7696_o;
  wire n7699_o;
  wire n7701_o;
  wire n7703_o;
  wire n7706_o;
  wire n7709_o;
  wire n7712_o;
  wire n7715_o;
  wire n7718_o;
  wire n7721_o;
  wire n7724_o;
  wire n7727_o;
  wire n7730_o;
  wire [1:0] n7732_o;
  wire [5:0] n7733_o;
  wire [5:0] n7734_o;
  wire n7736_o;
  wire n7738_o;
  wire n7740_o;
  wire n7744_o;
  wire n7747_o;
  wire n7750_o;
  wire n7753_o;
  wire n7756_o;
  wire n7759_o;
  wire n7762_o;
  wire n7765_o;
  wire n7768_o;
  wire n7771_o;
  wire n7774_o;
  wire n7777_o;
  wire [4:0] n7779_o;
  wire [2:0] n7780_o;
  wire [15:0] n7781_o;
  wire [1:0] n7782_o;
  wire [2:0] n7783_o;
  wire n7784_o;
  wire n7785_o;
  wire [2:0] n7786_o;
  wire [2:0] n7787_o;
  wire n7788_o;
  wire n7789_o;
  wire n7790_o;
  wire n7791_o;
  wire n7792_o;
  wire n7793_o;
  wire n7794_o;
  wire n7795_o;
  wire [1:0] n7796_o;
  wire [4:0] n7797_o;
  wire [2:0] n7799_o;
  wire [2:0] n7800_o;
  wire [15:0] n7801_o;
  wire [3:0] n7803_o;
  wire n7805_o;
  wire n7806_o;
  wire n7807_o;
  wire n7808_o;
  wire n7809_o;
  wire [1:0] n7810_o;
  wire n7812_o;
  wire n7813_o;
  wire n7814_o;
  wire n7815_o;
  wire [15:0] n7820_o;
  wire n7821_o;
  wire [3:0] n7826_o;
  wire n7827_o;
  wire n7828_o;
  wire n7831_o;
  wire n7832_o;
  wire n7836_o;
  wire [16:0] n7838_o;
  wire [4:0] n7839_o;
  wire [3:0] n7840_o;
  wire [16:0] n7842_o;
  wire n7844_o;
  wire n7846_o;
  localparam [4:0] n7847_o = 5'b00000;
  wire [3:0] n7850_o;
  wire n7852_o;
  localparam [88:0] n7853_o = 89'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  wire n7858_o;
  wire n7860_o;
  wire [39:0] n7862_o;
  wire [8:0] n7863_o;
  wire [6:0] n7864_o;
  wire n7865_o;
  wire n7866_o;
  wire n7867_o;
  wire n7868_o;
  wire [1:0] n7869_o;
  wire n7871_o;
  wire n7872_o;
  wire n7873_o;
  wire n7875_o;
  wire n7876_o;
  wire n7877_o;
  wire n7878_o;
  wire n7879_o;
  wire n7881_o;
  wire n7883_o;
  wire n7885_o;
  wire n7887_o;
  wire n7888_o;
  wire n7890_o;
  wire n7891_o;
  wire n7892_o;
  wire n7893_o;
  wire n7894_o;
  wire n7895_o;
  wire n7896_o;
  wire n7898_o;
  wire n7899_o;
  wire n7900_o;
  wire n7901_o;
  wire n7902_o;
  wire n7903_o;
  wire [3:0] n7904_o;
  wire [3:0] n7905_o;
  wire [3:0] n7906_o;
  wire n7909_o;
  wire [2:0] n7910_o;
  wire n7912_o;
  wire n7914_o;
  wire n7915_o;
  wire n7916_o;
  wire n7917_o;
  wire [1:0] n7921_o;
  wire n7923_o;
  wire n7924_o;
  wire n7925_o;
  wire n7926_o;
  wire n7927_o;
  wire n7928_o;
  wire n7929_o;
  wire n7930_o;
  wire n7931_o;
  wire n7932_o;
  wire n7933_o;
  wire n7934_o;
  wire n7935_o;
  wire [6:0] n7937_o;
  wire n7939_o;
  wire n7940_o;
  wire n7942_o;
  wire n7943_o;
  wire n7944_o;
  wire n7945_o;
  wire n7946_o;
  wire n7947_o;
  wire n7948_o;
  wire n7949_o;
  wire n7950_o;
  wire n7951_o;
  wire n7952_o;
  wire n7953_o;
  wire n7954_o;
  wire n7955_o;
  wire n7956_o;
  wire n7957_o;
  wire n7959_o;
  wire n7961_o;
  wire n7962_o;
  wire n7963_o;
  wire n7964_o;
  wire n7965_o;
  wire n7966_o;
  wire n7967_o;
  wire n7968_o;
  wire n7969_o;
  wire n7970_o;
  wire n7971_o;
  wire n7972_o;
  wire n7973_o;
  wire n7974_o;
  wire n7975_o;
  wire n7985_o;
  wire n7986_o;
  wire n7987_o;
  wire n7994_o;
  wire n7995_o;
  wire n7996_o;
  wire n7997_o;
  wire n7998_o;
  wire n8000_o;
  wire n8001_o;
  wire n8003_o;
  wire n8005_o;
  wire [6:0] n8006_o;
  wire n8007_o;
  wire [6:0] n8009_o;
  wire n8015_o;
  wire n8018_o;
  wire n8021_o;
  wire n8022_o;
  wire n8023_o;
  wire n8025_o;
  wire n8026_o;
  wire n8027_o;
  wire n8029_o;
  wire n8030_o;
  wire n8032_o;
  wire n8033_o;
  wire n8035_o;
  wire n8037_o;
  wire n8038_o;
  wire n8039_o;
  wire n8040_o;
  wire n8041_o;
  wire n8043_o;
  wire n8044_o;
  wire n8045_o;
  wire n8046_o;
  wire [1:0] n8048_o;
  wire n8049_o;
  wire n8050_o;
  wire n8051_o;
  wire n8052_o;
  wire [1:0] n8054_o;
  wire n8057_o;
  wire n8060_o;
  wire n8061_o;
  wire n8062_o;
  wire n8063_o;
  wire n8064_o;
  wire n8065_o;
  wire n8066_o;
  wire n8067_o;
  wire [6:0] n8070_o;
  wire n8072_o;
  wire n8075_o;
  wire n8076_o;
  wire n8079_o;
  wire n8080_o;
  wire n8081_o;
  wire n8082_o;
  wire n8083_o;
  wire n8084_o;
  wire [1:0] n8086_o;
  wire n8088_o;
  wire [6:0] n8091_o;
  wire [1:0] n8092_o;
  wire n8094_o;
  wire [1:0] n8098_o;
  wire n8101_o;
  wire n8103_o;
  wire n8104_o;
  wire n8105_o;
  wire n8106_o;
  wire n8107_o;
  wire n8108_o;
  wire [6:0] n8110_o;
  wire [1:0] n8112_o;
  wire n8114_o;
  wire n8115_o;
  wire n8116_o;
  wire n8117_o;
  wire n8118_o;
  wire n8119_o;
  wire n8120_o;
  wire n8121_o;
  wire [6:0] n8122_o;
  wire n8124_o;
  wire n8127_o;
  wire n8129_o;
  wire n8130_o;
  wire n8131_o;
  wire n8133_o;
  wire n8134_o;
  wire n8135_o;
  wire n8136_o;
  wire [1:0] n8138_o;
  wire n8139_o;
  wire n8140_o;
  wire n8141_o;
  wire n8142_o;
  wire n8144_o;
  wire n8145_o;
  wire n8148_o;
  wire n8149_o;
  wire n8150_o;
  wire n8151_o;
  wire n8152_o;
  wire [1:0] n8156_o;
  wire n8158_o;
  wire n8159_o;
  wire n8160_o;
  wire [6:0] n8162_o;
  wire n8164_o;
  wire n8166_o;
  wire n8167_o;
  wire n8168_o;
  wire n8170_o;
  wire n8171_o;
  wire n8172_o;
  wire n8174_o;
  wire n8175_o;
  wire n8177_o;
  wire n8179_o;
  wire n8180_o;
  wire n8181_o;
  wire n8182_o;
  wire n8184_o;
  wire n8185_o;
  wire n8186_o;
  wire n8187_o;
  wire [1:0] n8189_o;
  wire n8190_o;
  wire n8191_o;
  wire n8192_o;
  wire n8193_o;
  wire [1:0] n8195_o;
  wire n8198_o;
  wire n8201_o;
  wire n8202_o;
  wire n8203_o;
  wire n8204_o;
  wire n8205_o;
  wire n8206_o;
  wire n8207_o;
  wire [6:0] n8210_o;
  wire n8212_o;
  wire n8215_o;
  wire n8216_o;
  wire n8219_o;
  wire n8220_o;
  wire n8221_o;
  wire n8222_o;
  wire n8223_o;
  wire n8224_o;
  wire [1:0] n8226_o;
  wire n8228_o;
  wire [6:0] n8231_o;
  wire [1:0] n8232_o;
  wire n8234_o;
  wire [1:0] n8239_o;
  wire n8240_o;
  wire n8241_o;
  wire n8242_o;
  wire n8243_o;
  wire n8244_o;
  wire n8245_o;
  wire n8246_o;
  wire n8247_o;
  wire [6:0] n8250_o;
  wire [1:0] n8252_o;
  wire n8253_o;
  wire n8254_o;
  wire n8255_o;
  wire n8256_o;
  wire n8257_o;
  wire n8258_o;
  wire n8259_o;
  wire n8260_o;
  wire n8261_o;
  wire [6:0] n8262_o;
  wire n8264_o;
  wire n8268_o;
  wire n8271_o;
  wire n8272_o;
  wire n8273_o;
  wire n8275_o;
  wire n8276_o;
  wire n8277_o;
  wire n8278_o;
  wire [1:0] n8280_o;
  wire n8281_o;
  wire n8282_o;
  wire n8283_o;
  wire n8284_o;
  wire n8286_o;
  wire n8288_o;
  wire n8291_o;
  wire n8292_o;
  wire n8293_o;
  wire n8294_o;
  wire n8295_o;
  wire [1:0] n8299_o;
  wire n8300_o;
  wire [6:0] n8303_o;
  wire n8305_o;
  wire n8307_o;
  wire n8310_o;
  wire [6:0] n8312_o;
  wire n8314_o;
  wire n8316_o;
  wire n8317_o;
  wire n8320_o;
  wire n8323_o;
  wire n8325_o;
  wire n8326_o;
  wire n8327_o;
  wire n8329_o;
  wire n8332_o;
  wire [6:0] n8334_o;
  wire n8335_o;
  wire n8338_o;
  wire n8340_o;
  wire n8341_o;
  wire n8343_o;
  wire n8349_o;
  wire n8350_o;
  wire [1:0] n8351_o;
  wire n8353_o;
  wire n8355_o;
  wire n8356_o;
  wire [1:0] n8358_o;
  wire n8361_o;
  wire n8363_o;
  wire n8368_o;
  wire n8370_o;
  wire [1:0] n8372_o;
  wire n8375_o;
  wire n8379_o;
  wire n8380_o;
  wire [1:0] n8382_o;
  wire [6:0] n8384_o;
  wire n8386_o;
  wire n8388_o;
  wire n8389_o;
  wire n8391_o;
  wire n8393_o;
  wire n8395_o;
  wire n8396_o;
  wire [1:0] n8403_o;
  wire n8406_o;
  wire n8407_o;
  wire n8408_o;
  wire n8409_o;
  wire n8410_o;
  wire n8411_o;
  wire n8412_o;
  wire n8413_o;
  wire n8414_o;
  wire n8415_o;
  wire n8416_o;
  wire n8417_o;
  wire n8418_o;
  wire [6:0] n8420_o;
  wire n8422_o;
  wire n8423_o;
  wire n8426_o;
  wire n8432_o;
  wire n8435_o;
  wire n8436_o;
  wire n8438_o;
  wire n8439_o;
  wire n8440_o;
  wire n8441_o;
  wire n8447_o;
  wire n8450_o;
  wire n8451_o;
  wire n8453_o;
  wire [1:0] n8461_o;
  wire n8464_o;
  wire n8466_o;
  wire n8469_o;
  wire n8471_o;
  wire n8472_o;
  wire n8473_o;
  wire n8474_o;
  wire n8475_o;
  wire n8476_o;
  wire n8477_o;
  wire n8478_o;
  wire n8479_o;
  wire n8480_o;
  wire n8481_o;
  wire n8482_o;
  wire n8483_o;
  wire n8484_o;
  wire n8485_o;
  wire n8486_o;
  wire n8487_o;
  wire n8488_o;
  wire [6:0] n8491_o;
  wire n8493_o;
  wire n8497_o;
  wire n8501_o;
  wire [15:0] n8502_o;
  wire n8504_o;
  wire [2:0] n8505_o;
  wire n8507_o;
  wire n8509_o;
  wire n8511_o;
  wire n8512_o;
  wire n8513_o;
  wire n8514_o;
  wire n8515_o;
  wire n8516_o;
  wire [1:0] n8518_o;
  wire n8519_o;
  wire n8520_o;
  wire n8521_o;
  wire n8522_o;
  wire n8523_o;
  wire [6:0] n8525_o;
  wire n8527_o;
  wire n8528_o;
  wire n8531_o;
  wire n8532_o;
  wire [1:0] n8536_o;
  wire n8537_o;
  wire n8538_o;
  wire n8539_o;
  wire n8540_o;
  wire [1:0] n8542_o;
  wire n8543_o;
  wire n8544_o;
  wire n8545_o;
  wire n8546_o;
  wire n8547_o;
  wire n8548_o;
  wire n8549_o;
  wire n8550_o;
  wire n8551_o;
  wire [6:0] n8553_o;
  wire n8555_o;
  wire [1:0] n8556_o;
  wire n8558_o;
  wire n8560_o;
  wire n8562_o;
  wire [2:0] n8563_o;
  wire n8565_o;
  wire n8567_o;
  wire n8572_o;
  wire [2:0] n8573_o;
  wire n8575_o;
  wire n8577_o;
  wire [1:0] n8579_o;
  wire n8581_o;
  wire [1:0] n8584_o;
  wire n8587_o;
  wire n8589_o;
  wire [2:0] n8590_o;
  wire n8592_o;
  wire n8594_o;
  wire n8597_o;
  wire [2:0] n8598_o;
  wire n8600_o;
  wire n8602_o;
  wire n8605_o;
  wire n8609_o;
  wire n8612_o;
  wire n8615_o;
  wire n8618_o;
  wire n8621_o;
  wire n8624_o;
  wire n8625_o;
  wire n8627_o;
  wire [1:0] n8630_o;
  wire n8631_o;
  wire n8632_o;
  wire [6:0] n8635_o;
  wire n8637_o;
  wire n8638_o;
  wire n8640_o;
  wire n8643_o;
  wire n8646_o;
  wire n8650_o;
  wire n8653_o;
  wire n8656_o;
  wire n8659_o;
  wire n8662_o;
  wire n8665_o;
  wire n8668_o;
  wire n8671_o;
  wire n8674_o;
  wire n8675_o;
  wire n8676_o;
  wire n8679_o;
  wire n8680_o;
  wire n8681_o;
  wire n8682_o;
  wire n8683_o;
  wire n8685_o;
  wire n8687_o;
  wire n8688_o;
  wire n8689_o;
  wire [1:0] n8692_o;
  wire n8694_o;
  wire n8695_o;
  wire [6:0] n8698_o;
  wire n8700_o;
  wire n8702_o;
  wire [3:0] n8703_o;
  wire n8705_o;
  wire [1:0] n8709_o;
  wire [1:0] n8711_o;
  wire n8713_o;
  wire n8714_o;
  wire [6:0] n8717_o;
  wire n8719_o;
  wire n8721_o;
  wire n8723_o;
  wire n8726_o;
  wire [11:0] n8728_o;
  wire n8730_o;
  wire [11:0] n8731_o;
  wire n8733_o;
  wire n8734_o;
  wire [11:0] n8735_o;
  wire n8737_o;
  wire n8738_o;
  wire [11:0] n8739_o;
  wire n8741_o;
  wire n8742_o;
  wire n8743_o;
  wire [11:0] n8744_o;
  wire n8746_o;
  wire [11:0] n8747_o;
  wire n8749_o;
  wire n8750_o;
  wire [11:0] n8751_o;
  wire n8753_o;
  wire n8754_o;
  wire [11:0] n8755_o;
  wire n8757_o;
  wire n8758_o;
  wire n8759_o;
  wire n8760_o;
  wire n8761_o;
  wire n8762_o;
  wire n8764_o;
  wire n8766_o;
  wire n8768_o;
  wire n8769_o;
  wire n8771_o;
  wire n8775_o;
  wire n8777_o;
  wire n8778_o;
  wire n8779_o;
  wire n8780_o;
  wire n8781_o;
  wire n8782_o;
  wire [1:0] n8785_o;
  wire n8787_o;
  wire n8788_o;
  wire n8791_o;
  wire n8792_o;
  wire n8793_o;
  wire n8794_o;
  wire n8795_o;
  wire n8796_o;
  wire n8797_o;
  wire n8798_o;
  wire n8799_o;
  wire n8800_o;
  wire [1:0] n8803_o;
  wire n8805_o;
  wire n8806_o;
  wire n8810_o;
  wire n8811_o;
  wire [1:0] n8814_o;
  wire [1:0] n8816_o;
  wire [1:0] n8817_o;
  wire n8818_o;
  wire n8819_o;
  wire n8820_o;
  wire n8821_o;
  wire n8822_o;
  wire n8823_o;
  wire n8824_o;
  wire n8825_o;
  wire n8826_o;
  wire [6:0] n8828_o;
  wire n8830_o;
  wire n8831_o;
  wire n8832_o;
  wire [1:0] n8835_o;
  wire n8837_o;
  wire n8839_o;
  wire n8840_o;
  wire n8842_o;
  wire [5:0] n8845_o;
  wire n8847_o;
  wire n8850_o;
  wire [6:0] n8853_o;
  wire n8855_o;
  wire n8856_o;
  wire n8857_o;
  wire n8859_o;
  wire n8861_o;
  wire n8862_o;
  wire n8864_o;
  wire n8866_o;
  wire [1:0] n8868_o;
  wire [6:0] n8870_o;
  wire n8872_o;
  wire n8874_o;
  wire n8875_o;
  wire n8876_o;
  wire n8877_o;
  wire n8878_o;
  wire n8880_o;
  wire n8885_o;
  wire n8887_o;
  wire [15:0] n8888_o;
  wire n8890_o;
  wire n8891_o;
  wire n8892_o;
  wire n8894_o;
  wire [15:0] n8895_o;
  wire n8897_o;
  wire n8898_o;
  wire n8901_o;
  wire [6:0] n8903_o;
  wire n8906_o;
  wire n8907_o;
  wire n8909_o;
  wire [5:0] n8912_o;
  wire n8914_o;
  wire n8917_o;
  wire [6:0] n8920_o;
  wire n8922_o;
  wire n8923_o;
  wire n8924_o;
  wire n8925_o;
  wire n8927_o;
  wire n8928_o;
  wire n8929_o;
  wire n8931_o;
  wire [1:0] n8934_o;
  wire n8937_o;
  wire n8938_o;
  wire n8939_o;
  wire [6:0] n8941_o;
  wire n8944_o;
  wire n8945_o;
  wire n8948_o;
  wire n8949_o;
  wire n8950_o;
  wire n8951_o;
  wire n8952_o;
  wire n8955_o;
  wire [5:0] n8956_o;
  wire n8958_o;
  wire [5:0] n8959_o;
  wire [5:0] n8961_o;
  wire n8962_o;
  wire n8963_o;
  wire n8965_o;
  wire n8967_o;
  wire [84:0] n8968_o;
  reg n8971_o;
  reg [1:0] n8988_o;
  reg [1:0] n8989_o;
  reg [1:0] n9031_o;
  reg n9034_o;
  reg n9037_o;
  reg n9042_o;
  reg n9044_o;
  reg n9054_o;
  reg n9058_o;
  reg n9076_o;
  reg n9078_o;
  reg n9081_o;
  reg n9084_o;
  reg n9087_o;
  reg n9091_o;
  reg n9095_o;
  reg n9098_o;
  reg n9103_o;
  reg n9105_o;
  reg n9110_o;
  reg n9113_o;
  reg n9119_o;
  reg n9123_o;
  reg n9128_o;
  reg [5:0] n9129_o;
  reg n9133_o;
  reg n9136_o;
  reg n9140_o;
  reg n9142_o;
  reg n9143_o;
  reg n9146_o;
  reg n9148_o;
  reg n9150_o;
  wire n9151_o;
  reg n9152_o;
  wire n9153_o;
  reg n9154_o;
  reg n9155_o;
  reg n9156_o;
  reg n9157_o;
  reg n9158_o;
  wire n9159_o;
  reg n9160_o;
  reg n9161_o;
  reg n9162_o;
  wire n9163_o;
  wire n9164_o;
  wire n9165_o;
  reg n9166_o;
  reg n9167_o;
  wire n9168_o;
  wire n9169_o;
  wire n9170_o;
  reg n9171_o;
  wire n9172_o;
  wire n9173_o;
  wire n9174_o;
  reg n9175_o;
  reg n9176_o;
  reg n9177_o;
  reg n9178_o;
  wire n9179_o;
  wire n9180_o;
  wire n9181_o;
  reg n9182_o;
  reg n9183_o;
  wire n9184_o;
  wire n9185_o;
  wire n9186_o;
  reg n9187_o;
  wire n9188_o;
  wire n9189_o;
  wire n9190_o;
  reg n9191_o;
  wire n9192_o;
  wire n9193_o;
  wire n9194_o;
  reg n9195_o;
  wire n9196_o;
  wire n9197_o;
  wire n9198_o;
  reg n9199_o;
  reg n9200_o;
  wire n9201_o;
  wire n9202_o;
  wire n9203_o;
  reg n9204_o;
  wire n9205_o;
  reg n9206_o;
  wire n9207_o;
  reg n9208_o;
  reg n9209_o;
  reg n9210_o;
  reg n9211_o;
  wire n9212_o;
  wire n9213_o;
  wire n9214_o;
  reg n9215_o;
  wire n9216_o;
  reg n9217_o;
  reg n9218_o;
  reg n9219_o;
  wire n9220_o;
  wire n9221_o;
  wire n9222_o;
  reg n9223_o;
  wire n9224_o;
  wire n9225_o;
  wire n9226_o;
  reg n9227_o;
  wire n9228_o;
  wire n9229_o;
  wire n9230_o;
  reg n9231_o;
  wire n9232_o;
  reg n9233_o;
  wire n9234_o;
  reg n9235_o;
  wire n9237_o;
  wire n9238_o;
  wire n9239_o;
  wire n9240_o;
  wire n9244_o;
  wire n9245_o;
  wire n9246_o;
  wire [3:0] n9250_o;
  wire [3:0] n9251_o;
  wire [3:0] n9252_o;
  wire [2:0] n9259_o;
  wire [2:0] n9260_o;
  wire [2:0] n9261_o;
  wire [1:0] n9262_o;
  wire [1:0] n9263_o;
  wire [1:0] n9264_o;
  wire n9265_o;
  wire n9266_o;
  wire n9267_o;
  wire n9269_o;
  wire n9270_o;
  wire n9271_o;
  wire [3:0] n9272_o;
  wire n9280_o;
  reg n9281_o;
  wire [1:0] n9282_o;
  wire [5:0] n9283_o;
  reg [6:0] n9329_o;
  wire n9334_o;
  wire n9335_o;
  wire [11:0] n9336_o;
  wire [2:0] n9337_o;
  wire n9339_o;
  wire [2:0] n9340_o;
  wire n9342_o;
  wire [3:0] n9343_o;
  wire n9345_o;
  wire n9347_o;
  wire n9349_o;
  wire n9351_o;
  wire n9353_o;
  wire n9355_o;
  wire [7:0] n9356_o;
  reg [31:0] n9357_o;
  reg [3:0] n9358_o;
  reg [2:0] n9359_o;
  reg [2:0] n9360_o;
  wire [31:0] n9361_o;
  wire [3:0] n9362_o;
  wire [2:0] n9363_o;
  wire [2:0] n9364_o;
  wire [31:0] n9366_o;
  wire [3:0] n9368_o;
  wire [2:0] n9369_o;
  wire [2:0] n9370_o;
  wire [11:0] n9375_o;
  wire [31:0] n9377_o;
  wire n9379_o;
  wire [31:0] n9381_o;
  wire n9383_o;
  wire [3:0] n9385_o;
  wire [31:0] n9387_o;
  wire n9389_o;
  wire n9391_o;
  wire [3:0] n9392_o;
  reg [31:0] n9394_o;
  wire [3:0] n9399_o;
  wire n9401_o;
  wire n9403_o;
  wire n9404_o;
  wire n9405_o;
  wire n9406_o;
  wire n9407_o;
  wire n9408_o;
  wire n9410_o;
  wire n9411_o;
  wire n9412_o;
  wire n9413_o;
  wire n9415_o;
  wire n9416_o;
  wire n9417_o;
  wire n9419_o;
  wire n9420_o;
  wire n9422_o;
  wire n9423_o;
  wire n9424_o;
  wire n9426_o;
  wire n9427_o;
  wire n9429_o;
  wire n9430_o;
  wire n9431_o;
  wire n9433_o;
  wire n9434_o;
  wire n9436_o;
  wire n9437_o;
  wire n9438_o;
  wire n9440_o;
  wire n9441_o;
  wire n9443_o;
  wire n9444_o;
  wire n9445_o;
  wire n9446_o;
  wire n9447_o;
  wire n9448_o;
  wire n9449_o;
  wire n9450_o;
  wire n9451_o;
  wire n9452_o;
  wire n9454_o;
  wire n9455_o;
  wire n9456_o;
  wire n9457_o;
  wire n9458_o;
  wire n9459_o;
  wire n9460_o;
  wire n9461_o;
  wire n9462_o;
  wire n9463_o;
  wire n9465_o;
  wire n9466_o;
  wire n9467_o;
  wire n9468_o;
  wire n9469_o;
  wire n9470_o;
  wire n9471_o;
  wire n9472_o;
  wire n9473_o;
  wire n9474_o;
  wire n9475_o;
  wire n9476_o;
  wire n9477_o;
  wire n9478_o;
  wire n9479_o;
  wire n9480_o;
  wire n9482_o;
  wire n9483_o;
  wire n9484_o;
  wire n9485_o;
  wire n9486_o;
  wire n9487_o;
  wire n9488_o;
  wire n9489_o;
  wire n9490_o;
  wire n9491_o;
  wire n9492_o;
  wire n9493_o;
  wire n9495_o;
  wire [15:0] n9496_o;
  reg n9499_o;
  wire n9504_o;
  wire [15:0] n9505_o;
  wire n9506_o;
  wire n9507_o;
  wire n9508_o;
  wire n9511_o;
  wire n9514_o;
  wire n9517_o;
  wire n9520_o;
  wire n9523_o;
  wire n9526_o;
  wire n9529_o;
  wire n9532_o;
  wire n9535_o;
  wire n9538_o;
  wire n9541_o;
  wire n9544_o;
  wire n9547_o;
  wire n9550_o;
  wire n9553_o;
  wire n9556_o;
  wire [15:0] n9557_o;
  wire n9558_o;
  reg n9559_o;
  wire n9560_o;
  reg n9561_o;
  wire n9562_o;
  reg n9563_o;
  wire n9564_o;
  reg n9565_o;
  wire n9566_o;
  reg n9567_o;
  wire n9568_o;
  reg n9569_o;
  wire n9570_o;
  reg n9571_o;
  wire n9572_o;
  reg n9573_o;
  wire n9574_o;
  reg n9575_o;
  wire n9576_o;
  reg n9577_o;
  wire n9578_o;
  reg n9579_o;
  wire n9580_o;
  reg n9581_o;
  wire n9582_o;
  reg n9583_o;
  wire n9584_o;
  reg n9585_o;
  wire n9586_o;
  reg n9587_o;
  wire n9588_o;
  reg n9589_o;
  wire [15:0] n9590_o;
  wire [15:0] n9591_o;
  wire [15:0] n9592_o;
  wire [3:0] n9600_o;
  wire n9602_o;
  wire [3:0] n9603_o;
  wire n9605_o;
  wire [3:0] n9607_o;
  wire n9609_o;
  wire [3:0] n9610_o;
  wire n9612_o;
  wire n9615_o;
  wire [3:0] n9617_o;
  wire [3:0] n9618_o;
  wire n9620_o;
  wire [3:0] n9621_o;
  wire n9623_o;
  wire [3:0] n9624_o;
  wire [1:0] n9626_o;
  wire n9627_o;
  wire n9628_o;
  wire n9629_o;
  wire n9631_o;
  wire [3:0] n9632_o;
  wire n9634_o;
  wire [3:0] n9635_o;
  wire [1:0] n9636_o;
  wire [1:0] n9638_o;
  localparam [3:0] n9639_o = 4'b0000;
  wire [3:0] n9641_o;
  wire n9643_o;
  wire [1:0] n9645_o;
  wire n9647_o;
  wire n9649_o;
  wire n9650_o;
  wire n9652_o;
  wire n9653_o;
  wire n9654_o;
  wire n9655_o;
  wire n9657_o;
  wire n9658_o;
  wire [1:0] n9659_o;
  wire n9660_o;
  wire n9661_o;
  wire n9662_o;
  wire n9663_o;
  wire n9664_o;
  reg n9667_q;
  wire [3:0] n9668_o;
  reg [3:0] n9669_q;
  wire n9670_o;
  reg n9671_q;
  reg [31:0] n9672_q;
  wire [31:0] n9673_o;
  reg [31:0] n9674_q;
  wire [31:0] n9675_o;
  reg [31:0] n9676_q;
  reg [1:0] n9677_q;
  reg [1:0] n9678_q;
  reg n9679_q;
  reg [15:0] n9680_q;
  reg [15:0] n9681_q;
  wire [15:0] n9682_o;
  reg [15:0] n9683_q;
  reg [31:0] n9684_q;
  reg [31:0] n9685_q;
  reg [15:0] n9686_q;
  wire [3:0] n9688_o;
  reg [3:0] n9689_q;
  wire [31:0] n9690_o;
  wire [3:0] n9693_o;
  reg [3:0] n9694_q;
  wire [3:0] n9695_o;
  reg [3:0] n9696_q;
  wire n9697_o;
  reg n9698_q;
  wire [31:0] n9699_o;
  reg [31:0] n9700_q;
  wire [31:0] n9701_o;
  reg [31:0] n9702_q;
  wire n9703_o;
  reg n9704_q;
  reg [31:0] n9705_q;
  wire [31:0] n9706_o;
  reg [31:0] n9708_q;
  reg n9709_q;
  wire [31:0] n9711_o;
  reg n9712_q;
  reg [15:0] n9713_q;
  reg n9714_q;
  reg n9715_q;
  reg n9716_q;
  reg n9717_q;
  reg n9718_q;
  reg n9719_q;
  reg n9720_q;
  reg [7:0] n9721_q;
  reg n9722_q;
  wire n9723_o;
  reg n9724_q;
  reg [1:0] n9725_q;
  reg [5:0] n9726_q;
  wire n9727_o;
  reg n9728_q;
  wire [3:0] n9729_o;
  reg n9731_q;
  reg n9732_q;
  reg n9733_q;
  reg n9734_q;
  reg n9735_q;
  reg n9736_q;
  reg [7:0] n9737_q;
  reg n9738_q;
  reg n9739_q;
  reg n9740_q;
  reg n9741_q;
  wire [31:0] n9742_o;
  reg [31:0] n9743_q;
  wire [31:0] n9744_o;
  reg [31:0] n9745_q;
  reg [2:0] n9746_q;
  reg [7:0] n9747_q;
  reg n9748_q;
  reg n9749_q;
  reg n9750_q;
  reg n9751_q;
  reg n9752_q;
  wire [31:0] n9753_o;
  wire [7:0] n9754_o;
  reg [7:0] n9755_q;
  reg [5:0] n9756_q;
  reg [3:0] n9757_q;
  reg [5:0] n9758_q;
  reg n9759_q;
  reg n9760_q;
  reg [31:0] n9761_q;
  reg [31:0] n9762_q;
  wire [5:0] n9763_o;
  wire [5:0] n9764_o;
  reg [5:0] n9765_q;
  reg [5:0] n9766_q;
  wire [5:0] n9767_o;
  reg [31:0] n9768_q;
  reg [5:0] n9769_q;
  reg [31:0] n9770_q;
  reg [3:0] n9771_q;
  reg [2:0] n9772_q;
  reg [2:0] n9773_q;
  wire [88:0] n9774_o;
  wire [88:0] n9775_o;
  wire [88:0] n9776_o;
  reg [88:0] n9777_q;
  reg [6:0] n9778_q;
  reg n9779_q;
  reg [1:0] n9780_q;
  wire [2:0] n9781_o;
  wire [31:0] n9783_data; // mem_rd
  wire [31:0] n9784_data; // mem_rd
  assign addr_out = n1074_o;
  assign data_write = n278_o;
  assign nwr = n78_o;
  assign nuds = n89_o;
  assign nlds = n90_o;
  assign busstate = state;
  assign longword = n56_o;
  assign nresetout = n82_o;
  assign fc = n9781_o;
  assign clr_berr = n98_o;
  assign skipfetch = n8971_o;
  assign regin_out = regin;
  assign cacr_out = cacr;
  assign vbr_out = vbr;
  /* TG68KdotC_Kernel.vhd:148:16  */
  assign use_vbr_stackframe = n9667_q; // (signal)
  /* TG68KdotC_Kernel.vhd:150:16  */
  assign syncreset = n9669_q; // (signal)
  /* TG68KdotC_Kernel.vhd:151:16  */
  assign reset = n9671_q; // (signal)
  /* TG68KdotC_Kernel.vhd:152:16  */
  assign clkena_lw = n94_o; // (signal)
  /* TG68KdotC_Kernel.vhd:153:16  */
  assign tg68_pc = n9672_q; // (signal)
  /* TG68KdotC_Kernel.vhd:154:16  */
  assign tmp_tg68_pc = n9674_q; // (signal)
  /* TG68KdotC_Kernel.vhd:155:16  */
  assign tg68_pc_add = n1175_o; // (signal)
  /* TG68KdotC_Kernel.vhd:156:16  */
  assign pc_dataa = n1081_o; // (signal)
  /* TG68KdotC_Kernel.vhd:157:16  */
  assign pc_datab = n1174_o; // (signal)
  /* TG68KdotC_Kernel.vhd:158:16  */
  assign memaddr = n9676_q; // (signal)
  /* TG68KdotC_Kernel.vhd:159:16  */
  assign state = n9677_q; // (signal)
  /* TG68KdotC_Kernel.vhd:160:16  */
  assign datatype = n8988_o; // (signal)
  /* TG68KdotC_Kernel.vhd:161:16  */
  assign set_datatype = n8989_o; // (signal)
  /* TG68KdotC_Kernel.vhd:162:16  */
  assign exe_datatype = n9678_q; // (signal)
  /* TG68KdotC_Kernel.vhd:163:16  */
  assign setstate = n9031_o; // (signal)
  /* TG68KdotC_Kernel.vhd:164:16  */
  assign setaddrvalue = n9034_o; // (signal)
  /* TG68KdotC_Kernel.vhd:165:16  */
  assign addrvalue = n9679_q; // (signal)
  /* TG68KdotC_Kernel.vhd:167:16  */
  assign opcode = n9680_q; // (signal)
  /* TG68KdotC_Kernel.vhd:168:16  */
  assign exe_opcode = n9681_q; // (signal)
  /* TG68KdotC_Kernel.vhd:169:16  */
  assign sndopc = n9683_q; // (signal)
  /* TG68KdotC_Kernel.vhd:171:16  */
  assign exe_pc = n9684_q; // (signal)
  /* TG68KdotC_Kernel.vhd:172:16  */
  assign last_opc_pc = n9685_q; // (signal)
  /* TG68KdotC_Kernel.vhd:173:16  */
  assign last_opc_read = n9686_q; // (signal)
  /* TG68KdotC_Kernel.vhd:175:16  */
  assign reg_qa = n9784_data; // (signal)
  /* TG68KdotC_Kernel.vhd:176:16  */
  assign reg_qb = n9783_data; // (signal)
  /* TG68KdotC_Kernel.vhd:177:16  */
  assign wwrena = n392_o; // (signal)
  /* TG68KdotC_Kernel.vhd:177:23  */
  assign lwrena = n395_o; // (signal)
  /* TG68KdotC_Kernel.vhd:178:16  */
  assign bwrena = n398_o; // (signal)
  /* TG68KdotC_Kernel.vhd:179:16  */
  assign regwrena_now = n9037_o; // (signal)
  /* TG68KdotC_Kernel.vhd:180:16  */
  assign rf_dest_addr = n440_o; // (signal)
  /* TG68KdotC_Kernel.vhd:181:16  */
  assign rf_source_addr = n478_o; // (signal)
  /* TG68KdotC_Kernel.vhd:182:16  */
  assign rf_source_addrd = n9689_q; // (signal)
  /* TG68KdotC_Kernel.vhd:184:16  */
  assign regin = n9690_o; // (signal)
  /* TG68KdotC_Kernel.vhd:187:16  */
  assign rdindex_a = n9694_q; // (signal)
  /* TG68KdotC_Kernel.vhd:188:16  */
  assign rdindex_b = n9696_q; // (signal)
  /* TG68KdotC_Kernel.vhd:189:16  */
  assign wr_areg = n9698_q; // (signal)
  /* TG68KdotC_Kernel.vhd:192:16  */
  assign addr = n1073_o; // (signal)
  /* TG68KdotC_Kernel.vhd:193:16  */
  assign memaddr_reg = n1077_o; // (signal)
  /* TG68KdotC_Kernel.vhd:194:16  */
  assign memaddr_delta = n1072_o; // (signal)
  /* TG68KdotC_Kernel.vhd:195:16  */
  assign memaddr_delta_rega = n9700_q; // (signal)
  /* TG68KdotC_Kernel.vhd:196:16  */
  assign memaddr_delta_regb = n9702_q; // (signal)
  /* TG68KdotC_Kernel.vhd:197:16  */
  assign use_base = n9704_q; // (signal)
  /* TG68KdotC_Kernel.vhd:199:16  */
  assign ea_data = n9705_q; // (signal)
  /* TG68KdotC_Kernel.vhd:200:16  */
  assign op1out = n494_o; // (signal)
  /* TG68KdotC_Kernel.vhd:201:16  */
  assign op2out = n9706_o; // (signal)
  /* TG68KdotC_Kernel.vhd:202:16  */
  assign op1outbrief = n839_o; // (signal)
  /* TG68KdotC_Kernel.vhd:204:16  */
  assign aluout = alu_n42; // (signal)
  /* TG68KdotC_Kernel.vhd:205:16  */
  assign data_write_tmp = n9708_q; // (signal)
  /* TG68KdotC_Kernel.vhd:206:16  */
  assign data_write_muxin = n241_o; // (signal)
  /* TG68KdotC_Kernel.vhd:207:16  */
  assign data_write_mux = n250_o; // (signal)
  /* TG68KdotC_Kernel.vhd:208:16  */
  assign nextpass = n9709_q; // (signal)
  /* TG68KdotC_Kernel.vhd:209:16  */
  assign setnextpass = n9042_o; // (signal)
  /* TG68KdotC_Kernel.vhd:210:16  */
  assign setdispbyte = n9044_o; // (signal)
  /* TG68KdotC_Kernel.vhd:211:16  */
  assign setdisp = n9054_o; // (signal)
  /* TG68KdotC_Kernel.vhd:212:16  */
  assign regdirectsource = n7692_o; // (signal)
  /* TG68KdotC_Kernel.vhd:213:16  */
  assign addsub_q = alu_n41; // (signal)
  /* TG68KdotC_Kernel.vhd:214:16  */
  assign briefdata = n875_o; // (signal)
  /* TG68KdotC_Kernel.vhd:215:16  */
  assign c_out = alu_n40; // (signal)
  /* TG68KdotC_Kernel.vhd:218:16  */
  assign memaddr_a = n9711_o; // (signal)
  /* TG68KdotC_Kernel.vhd:220:16  */
  assign tg68_pc_brw = n9058_o; // (signal)
  /* TG68KdotC_Kernel.vhd:221:16  */
  assign tg68_pc_word = n9712_q; // (signal)
  /* TG68KdotC_Kernel.vhd:222:16  */
  assign getbrief = n7694_o; // (signal)
  /* TG68KdotC_Kernel.vhd:223:16  */
  assign brief = n9713_q; // (signal)
  /* TG68KdotC_Kernel.vhd:224:16  */
  assign data_is_source = n7696_o; // (signal)
  /* TG68KdotC_Kernel.vhd:225:16  */
  assign store_in_tmp = n9714_q; // (signal)
  /* TG68KdotC_Kernel.vhd:226:16  */
  assign write_back = n7959_o; // (signal)
  /* TG68KdotC_Kernel.vhd:227:16  */
  assign exec_write_back = n9715_q; // (signal)
  /* TG68KdotC_Kernel.vhd:228:16  */
  assign setstackaddr = n9076_o; // (signal)
  /* TG68KdotC_Kernel.vhd:229:16  */
  assign writepc = n9078_o; // (signal)
  /* TG68KdotC_Kernel.vhd:230:16  */
  assign writepcbig = n9716_q; // (signal)
  /* TG68KdotC_Kernel.vhd:231:16  */
  assign set_writepcbig = n9081_o; // (signal)
  /* TG68KdotC_Kernel.vhd:232:16  */
  assign writepcnext = n9717_q; // (signal)
  /* TG68KdotC_Kernel.vhd:233:16  */
  assign setopcode = n1211_o; // (signal)
  /* TG68KdotC_Kernel.vhd:234:16  */
  assign decodeopc = n9718_q; // (signal)
  /* TG68KdotC_Kernel.vhd:235:16  */
  assign execopc = n9719_q; // (signal)
  /* TG68KdotC_Kernel.vhd:236:16  */
  assign execopc_alu = n60_o; // (signal)
  /* TG68KdotC_Kernel.vhd:237:16  */
  assign setexecopc = n1236_o; // (signal)
  /* TG68KdotC_Kernel.vhd:238:16  */
  assign endopc = n9720_q; // (signal)
  /* TG68KdotC_Kernel.vhd:239:16  */
  assign setendopc = n1215_o; // (signal)
  /* TG68KdotC_Kernel.vhd:240:16  */
  assign flags = alu_n39; // (signal)
  /* TG68KdotC_Kernel.vhd:241:16  */
  assign flagssr = n9721_q; // (signal)
  /* TG68KdotC_Kernel.vhd:242:16  */
  assign srin = n1785_o; // (signal)
  /* TG68KdotC_Kernel.vhd:243:16  */
  assign exec_direct = n9722_q; // (signal)
  /* TG68KdotC_Kernel.vhd:244:16  */
  assign exec_tas = n9724_q; // (signal)
  /* TG68KdotC_Kernel.vhd:245:16  */
  assign set_exec_tas = n7706_o; // (signal)
  /* TG68KdotC_Kernel.vhd:247:16  */
  assign exe_condition = n9499_o; // (signal)
  /* TG68KdotC_Kernel.vhd:248:16  */
  assign ea_only = n7709_o; // (signal)
  /* TG68KdotC_Kernel.vhd:249:16  */
  assign source_areg = n9084_o; // (signal)
  /* TG68KdotC_Kernel.vhd:250:16  */
  assign source_lowbits = n7961_o; // (signal)
  /* TG68KdotC_Kernel.vhd:251:16  */
  assign source_ldrlbits = n9087_o; // (signal)
  /* TG68KdotC_Kernel.vhd:252:16  */
  assign source_ldrmbits = n9091_o; // (signal)
  /* TG68KdotC_Kernel.vhd:253:16  */
  assign source_2ndhbits = n7718_o; // (signal)
  /* TG68KdotC_Kernel.vhd:254:16  */
  assign source_2ndmbits = n9095_o; // (signal)
  /* TG68KdotC_Kernel.vhd:255:16  */
  assign source_2ndlbits = n9098_o; // (signal)
  /* TG68KdotC_Kernel.vhd:256:16  */
  assign dest_areg = n9103_o; // (signal)
  /* TG68KdotC_Kernel.vhd:257:16  */
  assign dest_ldrareg = n9105_o; // (signal)
  /* TG68KdotC_Kernel.vhd:258:16  */
  assign dest_ldrhbits = n9110_o; // (signal)
  /* TG68KdotC_Kernel.vhd:259:16  */
  assign dest_ldrlbits = n9113_o; // (signal)
  /* TG68KdotC_Kernel.vhd:260:16  */
  assign dest_2ndhbits = n9119_o; // (signal)
  /* TG68KdotC_Kernel.vhd:261:16  */
  assign dest_2ndlbits = n9123_o; // (signal)
  /* TG68KdotC_Kernel.vhd:262:16  */
  assign dest_hbits = n9128_o; // (signal)
  /* TG68KdotC_Kernel.vhd:263:16  */
  assign rot_bits = n9725_q; // (signal)
  /* TG68KdotC_Kernel.vhd:264:16  */
  assign set_rot_bits = n7732_o; // (signal)
  /* TG68KdotC_Kernel.vhd:265:16  */
  assign rot_cnt = n9726_q; // (signal)
  /* TG68KdotC_Kernel.vhd:266:16  */
  assign set_rot_cnt = n9129_o; // (signal)
  /* TG68KdotC_Kernel.vhd:267:16  */
  assign movem_actiond = n9728_q; // (signal)
  /* TG68KdotC_Kernel.vhd:268:16  */
  assign movem_regaddr = n9729_o; // (signal)
  /* TG68KdotC_Kernel.vhd:269:16  */
  assign movem_mux = n9641_o; // (signal)
  /* TG68KdotC_Kernel.vhd:270:16  */
  assign movem_presub = n7736_o; // (signal)
  /* TG68KdotC_Kernel.vhd:271:16  */
  assign movem_run = n9643_o; // (signal)
  /* TG68KdotC_Kernel.vhd:273:16  */
  assign set_direct_data = n9133_o; // (signal)
  /* TG68KdotC_Kernel.vhd:274:16  */
  assign use_direct_data = n9731_q; // (signal)
  /* TG68KdotC_Kernel.vhd:275:16  */
  assign direct_data = n9732_q; // (signal)
  /* TG68KdotC_Kernel.vhd:277:16  */
  assign set_v_flag = alu_n38; // (signal)
  /* TG68KdotC_Kernel.vhd:278:16  */
  assign set_vectoraddr = n9136_o; // (signal)
  /* TG68KdotC_Kernel.vhd:279:16  */
  assign writesr = n9140_o; // (signal)
  /* TG68KdotC_Kernel.vhd:280:16  */
  assign trap_berr = n9733_q; // (signal)
  /* TG68KdotC_Kernel.vhd:281:16  */
  assign trap_illegal = n9142_o; // (signal)
  /* TG68KdotC_Kernel.vhd:282:16  */
  assign trap_addr_error = n7744_o; // (signal)
  /* TG68KdotC_Kernel.vhd:283:16  */
  assign trap_priv = n7747_o; // (signal)
  /* TG68KdotC_Kernel.vhd:284:16  */
  assign trap_trace = n9734_q; // (signal)
  /* TG68KdotC_Kernel.vhd:285:16  */
  assign trap_1010 = n7750_o; // (signal)
  /* TG68KdotC_Kernel.vhd:286:16  */
  assign trap_1111 = n7753_o; // (signal)
  /* TG68KdotC_Kernel.vhd:287:16  */
  assign trap_trap = n7756_o; // (signal)
  /* TG68KdotC_Kernel.vhd:288:16  */
  assign trap_trapv = n7759_o; // (signal)
  /* TG68KdotC_Kernel.vhd:289:16  */
  assign trap_interrupt = n9735_q; // (signal)
  /* TG68KdotC_Kernel.vhd:290:16  */
  assign trapmake = n9143_o; // (signal)
  /* TG68KdotC_Kernel.vhd:291:16  */
  assign trapd = n9736_q; // (signal)
  /* TG68KdotC_Kernel.vhd:292:16  */
  assign trap_sr = n9737_q; // (signal)
  /* TG68KdotC_Kernel.vhd:293:16  */
  assign make_trace = n9738_q; // (signal)
  /* TG68KdotC_Kernel.vhd:294:16  */
  assign make_berr = n9739_q; // (signal)
  /* TG68KdotC_Kernel.vhd:295:16  */
  assign usestackframe2 = n9740_q; // (signal)
  /* TG68KdotC_Kernel.vhd:297:16  */
  assign set_stop = n7765_o; // (signal)
  /* TG68KdotC_Kernel.vhd:298:16  */
  assign stop = n9741_q; // (signal)
  /* TG68KdotC_Kernel.vhd:299:16  */
  assign trap_vector = n9743_q; // (signal)
  /* TG68KdotC_Kernel.vhd:300:16  */
  assign trap_vector_vbr = n917_o; // (signal)
  /* TG68KdotC_Kernel.vhd:301:16  */
  assign usp = n9745_q; // (signal)
  /* TG68KdotC_Kernel.vhd:306:16  */
  assign ipl_nr = n1238_o; // (signal)
  /* TG68KdotC_Kernel.vhd:307:16  */
  assign ripl_nr = n9746_q; // (signal)
  /* TG68KdotC_Kernel.vhd:308:16  */
  assign ipl_vec = n9747_q; // (signal)
  /* TG68KdotC_Kernel.vhd:309:16  */
  assign interrupt = n9748_q; // (signal)
  /* TG68KdotC_Kernel.vhd:310:16  */
  assign setinterrupt = n1218_o; // (signal)
  /* TG68KdotC_Kernel.vhd:311:16  */
  assign svmode = n9749_q; // (signal)
  /* TG68KdotC_Kernel.vhd:312:16  */
  assign presvmode = n9750_q; // (signal)
  /* TG68KdotC_Kernel.vhd:313:16  */
  assign suppress_base = n9751_q; // (signal)
  /* TG68KdotC_Kernel.vhd:314:16  */
  assign set_suppress_base = n9146_o; // (signal)
  /* TG68KdotC_Kernel.vhd:315:16  */
  assign set_z_error = n9148_o; // (signal)
  /* TG68KdotC_Kernel.vhd:316:16  */
  assign z_error = n9752_q; // (signal)
  /* TG68KdotC_Kernel.vhd:317:16  */
  assign ea_build_now = n7898_o; // (signal)
  /* TG68KdotC_Kernel.vhd:318:16  */
  assign build_logical = n7771_o; // (signal)
  /* TG68KdotC_Kernel.vhd:319:16  */
  assign build_bcd = n7774_o; // (signal)
  /* TG68KdotC_Kernel.vhd:321:16  */
  assign data_read = n9753_o; // (signal)
  /* TG68KdotC_Kernel.vhd:322:16  */
  assign bf_ext_in = n9755_q; // (signal)
  /* TG68KdotC_Kernel.vhd:323:16  */
  assign bf_ext_out = alu_n36; // (signal)
  /* TG68KdotC_Kernel.vhd:325:16  */
  assign long_start = n234_o; // (signal)
  /* TG68KdotC_Kernel.vhd:326:16  */
  assign long_start_alu = n58_o; // (signal)
  /* TG68KdotC_Kernel.vhd:327:16  */
  assign non_aligned = n72_o; // (signal)
  /* TG68KdotC_Kernel.vhd:328:16  */
  assign check_aligned = n7777_o; // (signal)
  /* TG68KdotC_Kernel.vhd:329:16  */
  assign long_done = n236_o; // (signal)
  /* TG68KdotC_Kernel.vhd:330:16  */
  assign memmask = n9756_q; // (signal)
  /* TG68KdotC_Kernel.vhd:331:16  */
  assign set_memmask = n1769_o; // (signal)
  /* TG68KdotC_Kernel.vhd:332:16  */
  assign memread = n9757_q; // (signal)
  /* TG68KdotC_Kernel.vhd:333:16  */
  assign wbmemmask = n9758_q; // (signal)
  /* TG68KdotC_Kernel.vhd:334:16  */
  assign memmaskmux = n85_o; // (signal)
  /* TG68KdotC_Kernel.vhd:335:16  */
  assign oddout = n9759_q; // (signal)
  /* TG68KdotC_Kernel.vhd:336:16  */
  assign set_oddout = n1694_o; // (signal)
  /* TG68KdotC_Kernel.vhd:337:16  */
  assign pcbase = n9760_q; // (signal)
  /* TG68KdotC_Kernel.vhd:338:16  */
  assign set_pcbase = n2160_o; // (signal)
  /* TG68KdotC_Kernel.vhd:340:16  */
  assign last_data_read = n9761_q; // (signal)
  /* TG68KdotC_Kernel.vhd:341:16  */
  assign last_data_in = n9762_q; // (signal)
  /* TG68KdotC_Kernel.vhd:343:16  */
  assign bf_offset = n9763_o; // (signal)
  /* TG68KdotC_Kernel.vhd:344:16  */
  assign bf_width = n9764_o; // (signal)
  /* TG68KdotC_Kernel.vhd:345:16  */
  assign bf_bhits = n1692_o; // (signal)
  /* TG68KdotC_Kernel.vhd:346:16  */
  assign bf_shift = n1749_o; // (signal)
  /* TG68KdotC_Kernel.vhd:347:16  */
  assign alu_width = n9765_q; // (signal)
  /* TG68KdotC_Kernel.vhd:348:16  */
  assign alu_bf_shift = n9766_q; // (signal)
  /* TG68KdotC_Kernel.vhd:349:16  */
  assign bf_loffset = n9767_o; // (signal)
  /* TG68KdotC_Kernel.vhd:350:16  */
  assign bf_full_offset = n1682_o; // (signal)
  /* TG68KdotC_Kernel.vhd:351:16  */
  assign alu_bf_ffo_offset = n9768_q; // (signal)
  /* TG68KdotC_Kernel.vhd:352:16  */
  assign alu_bf_loffset = n9769_q; // (signal)
  /* TG68KdotC_Kernel.vhd:354:16  */
  assign movec_data = n9394_o; // (signal)
  /* TG68KdotC_Kernel.vhd:355:16  */
  assign vbr = n9770_q; // (signal)
  /* TG68KdotC_Kernel.vhd:356:16  */
  assign cacr = n9771_q; // (signal)
  /* TG68KdotC_Kernel.vhd:357:16  */
  assign dfc = n9772_q; // (signal)
  /* TG68KdotC_Kernel.vhd:358:16  */
  assign sfc = n9773_q; // (signal)
  /* TG68KdotC_Kernel.vhd:361:16  */
  assign set = n9774_o; // (signal)
  /* TG68KdotC_Kernel.vhd:362:16  */
  assign set_exec = n9775_o; // (signal)
  /* TG68KdotC_Kernel.vhd:363:16  */
  assign exec = n9777_q; // (signal)
  /* TG68KdotC_Kernel.vhd:365:16  */
  assign micro_state = n9778_q; // (signal)
  /* TG68KdotC_Kernel.vhd:366:16  */
  assign next_micro_state = n9329_o; // (signal)
  /* TG68KdotC_Kernel.vhd:405:49  */
  assign n34_o = last_data_read[15:0];
  /* TG68KdotC_Kernel.vhd:406:39  */
  assign n35_o = data_read[15:0];
  /* TG68KdotC_Kernel.vhd:410:31  */
  assign alu_n36 = alu_bf_ext_out; // (signal)
  /* TG68KdotC_Kernel.vhd:414:45  */
  assign n37_o = alu_bf_loffset[4:0];
  /* TG68KdotC_Kernel.vhd:416:31  */
  assign alu_n38 = alu_set_v_flag; // (signal)
  /* TG68KdotC_Kernel.vhd:417:26  */
  assign alu_n39 = alu_flags; // (signal)
  /* TG68KdotC_Kernel.vhd:418:26  */
  assign alu_n40 = alu_c_out; // (signal)
  /* TG68KdotC_Kernel.vhd:419:29  */
  assign alu_n41 = alu_addsub_q; // (signal)
  /* TG68KdotC_Kernel.vhd:420:27  */
  assign alu_n42 = alu_aluout; // (signal)
  /* TG68KdotC_Kernel.vhd:372:1  */
  tg68k_alu_2_0_2_0 alu (
    .clk(clk),
    .reset(reset),
    .clkena_lw(clkena_lw),
    .cpu(cpu),
    .execopc(execopc_alu),
    .decodeopc(decodeopc),
    .exe_condition(exe_condition),
    .exec_tas(exec_tas),
    .long_start(long_start_alu),
    .non_aligned(non_aligned),
    .check_aligned(check_aligned),
    .movem_presub(movem_presub),
    .set_stop(set_stop),
    .z_error(z_error),
    .rot_bits(rot_bits),
    .exec(exec),
    .op1out(op1out),
    .op2out(op2out),
    .reg_qa(reg_qa),
    .reg_qb(reg_qb),
    .opcode(opcode),
    .exe_opcode(exe_opcode),
    .exe_datatype(exe_datatype),
    .sndopc(sndopc),
    .last_data_read(n34_o),
    .data_read(n35_o),
    .flagssr(flagssr),
    .micro_state(micro_state),
    .bf_ext_in(bf_ext_in),
    .bf_shift(alu_bf_shift),
    .bf_width(alu_width),
    .bf_ffo_offset(alu_bf_ffo_offset),
    .bf_loffset(n37_o),
    .bf_ext_out(alu_bf_ext_out),
    .set_v_flag(alu_set_v_flag),
    .flags(alu_flags),
    .c_out(alu_c_out),
    .addsub_q(alu_addsub_q),
    .aluout(alu_aluout));
  /* TG68KdotC_Kernel.vhd:424:35  */
  assign n55_o = memmaskmux[3];
  /* TG68KdotC_Kernel.vhd:424:21  */
  assign n56_o = ~n55_o;
  /* TG68KdotC_Kernel.vhd:426:48  */
  assign n57_o = memmaskmux[3];
  /* TG68KdotC_Kernel.vhd:426:34  */
  assign n58_o = ~n57_o;
  /* TG68KdotC_Kernel.vhd:427:39  */
  assign n59_o = exec[84];
  /* TG68KdotC_Kernel.vhd:427:32  */
  assign n60_o = execopc | n59_o;
  /* TG68KdotC_Kernel.vhd:431:31  */
  assign n63_o = memmaskmux[5:4];
  /* TG68KdotC_Kernel.vhd:431:44  */
  assign n65_o = n63_o == 2'b01;
  /* TG68KdotC_Kernel.vhd:431:66  */
  assign n66_o = memmaskmux[5:4];
  /* TG68KdotC_Kernel.vhd:431:79  */
  assign n68_o = n66_o == 2'b10;
  /* TG68KdotC_Kernel.vhd:431:52  */
  assign n69_o = n65_o | n68_o;
  /* TG68KdotC_Kernel.vhd:431:17  */
  assign n72_o = n69_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:441:30  */
  assign n77_o = state == 2'b11;
  /* TG68KdotC_Kernel.vhd:441:20  */
  assign n78_o = n77_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:443:35  */
  assign n81_o = exec[74];
  /* TG68KdotC_Kernel.vhd:443:26  */
  assign n82_o = n81_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:447:40  */
  assign n84_o = addr[0];
  /* TG68KdotC_Kernel.vhd:447:31  */
  assign n85_o = n84_o ? memmask : n88_o;
  /* TG68KdotC_Kernel.vhd:447:62  */
  assign n86_o = memmask[4:0];
  /* TG68KdotC_Kernel.vhd:447:75  */
  assign n88_o = {n86_o, 1'b1};
  /* TG68KdotC_Kernel.vhd:448:27  */
  assign n89_o = memmaskmux[5];
  /* TG68KdotC_Kernel.vhd:449:27  */
  assign n90_o = memmaskmux[4];
  /* TG68KdotC_Kernel.vhd:450:59  */
  assign n92_o = memmaskmux[3];
  /* TG68KdotC_Kernel.vhd:450:45  */
  assign n93_o = n92_o & clkena_in;
  /* TG68KdotC_Kernel.vhd:450:26  */
  assign n94_o = n93_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:451:44  */
  assign n97_o = trap_berr & setopcode;
  /* TG68KdotC_Kernel.vhd:451:25  */
  assign n98_o = n97_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:455:26  */
  assign n102_o = ~nreset;
  /* TG68KdotC_Kernel.vhd:460:55  */
  assign n104_o = syncreset[2:0];
  /* TG68KdotC_Kernel.vhd:460:67  */
  assign n106_o = {n104_o, 1'b1};
  /* TG68KdotC_Kernel.vhd:461:55  */
  assign n107_o = syncreset[3];
  /* TG68KdotC_Kernel.vhd:461:42  */
  assign n108_o = ~n107_o;
  /* TG68KdotC_Kernel.vhd:465:52  */
  assign n118_o = cpu[0];
  /* TG68KdotC_Kernel.vhd:465:60  */
  assign n120_o = 1'b1 & n118_o;
  /* TG68KdotC_Kernel.vhd:465:45  */
  assign n122_o = 1'b0 | n120_o;
  /* TG68KdotC_Kernel.vhd:465:25  */
  assign n125_o = n122_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:475:30  */
  assign n130_o = memmaskmux[4];
  /* TG68KdotC_Kernel.vhd:475:33  */
  assign n131_o = ~n130_o;
  /* TG68KdotC_Kernel.vhd:476:50  */
  assign n132_o = last_data_in[15:0];
  /* TG68KdotC_Kernel.vhd:476:63  */
  assign n133_o = {n132_o, data_in};
  /* TG68KdotC_Kernel.vhd:478:50  */
  assign n134_o = last_data_in[23:0];
  /* TG68KdotC_Kernel.vhd:478:71  */
  assign n135_o = data_in[15:8];
  /* TG68KdotC_Kernel.vhd:478:63  */
  assign n136_o = {n134_o, n135_o};
  /* TG68KdotC_Kernel.vhd:480:27  */
  assign n138_o = memread[0];
  /* TG68KdotC_Kernel.vhd:480:46  */
  assign n139_o = memread[1:0];
  /* TG68KdotC_Kernel.vhd:480:58  */
  assign n141_o = n139_o == 2'b10;
  /* TG68KdotC_Kernel.vhd:480:78  */
  assign n142_o = memmaskmux[4];
  /* TG68KdotC_Kernel.vhd:480:64  */
  assign n143_o = n142_o & n141_o;
  /* TG68KdotC_Kernel.vhd:480:35  */
  assign n144_o = n138_o | n143_o;
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n145_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n146_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n147_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n148_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n149_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n150_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n151_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n152_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n153_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n154_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n155_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n156_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n157_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n158_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n159_o = data_read[15];
  /* TG68KdotC_Kernel.vhd:481:70  */
  assign n160_o = data_read[15];
  assign n161_o = {n145_o, n146_o, n147_o, n148_o};
  assign n162_o = {n149_o, n150_o, n151_o, n152_o};
  assign n163_o = {n153_o, n154_o, n155_o, n156_o};
  assign n164_o = {n157_o, n158_o, n159_o, n160_o};
  assign n165_o = {n161_o, n162_o, n163_o, n164_o};
  assign n166_o = n133_o[31:16];
  assign n167_o = n136_o[31:16];
  /* TG68KdotC_Kernel.vhd:475:17  */
  assign n168_o = n131_o ? n166_o : n167_o;
  /* TG68KdotC_Kernel.vhd:480:17  */
  assign n169_o = n144_o ? n165_o : n168_o;
  assign n170_o = n133_o[15:0];
  assign n171_o = n136_o[15:0];
  /* TG68KdotC_Kernel.vhd:475:17  */
  assign n172_o = n131_o ? n170_o : n171_o;
  /* TG68KdotC_Kernel.vhd:485:51  */
  assign n175_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:485:42  */
  assign n176_o = n175_o & clkena_lw;
  /* TG68KdotC_Kernel.vhd:486:46  */
  assign n177_o = memmaskmux[4];
  /* TG68KdotC_Kernel.vhd:486:49  */
  assign n178_o = ~n177_o;
  /* TG68KdotC_Kernel.vhd:487:66  */
  assign n179_o = last_data_in[23:16];
  /* TG68KdotC_Kernel.vhd:489:66  */
  assign n180_o = last_data_in[31:24];
  /* TG68KdotC_Kernel.vhd:486:33  */
  assign n181_o = n178_o ? n179_o : n180_o;
  /* TG68KdotC_Kernel.vhd:495:41  */
  assign n184_o = state == 2'b00;
  /* TG68KdotC_Kernel.vhd:495:54  */
  assign n185_o = exec[38];
  /* TG68KdotC_Kernel.vhd:495:47  */
  assign n186_o = n184_o | n185_o;
  /* TG68KdotC_Kernel.vhd:497:49  */
  assign n187_o = state[1];
  /* TG68KdotC_Kernel.vhd:497:52  */
  assign n188_o = ~n187_o;
  /* TG68KdotC_Kernel.vhd:497:68  */
  assign n189_o = memmask[1];
  /* TG68KdotC_Kernel.vhd:497:71  */
  assign n190_o = ~n189_o;
  /* TG68KdotC_Kernel.vhd:497:57  */
  assign n191_o = n190_o & n188_o;
  /* TG68KdotC_Kernel.vhd:499:52  */
  assign n192_o = state[1];
  /* TG68KdotC_Kernel.vhd:499:55  */
  assign n193_o = ~n192_o;
  /* TG68KdotC_Kernel.vhd:499:70  */
  assign n194_o = memread[1];
  /* TG68KdotC_Kernel.vhd:499:60  */
  assign n195_o = n193_o | n194_o;
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n196_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n197_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n198_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n199_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n200_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n201_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n202_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n203_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n204_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n205_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n206_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n207_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n208_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n209_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n210_o = data_in[15];
  /* TG68KdotC_Kernel.vhd:500:97  */
  assign n211_o = data_in[15];
  assign n212_o = {n196_o, n197_o, n198_o, n199_o};
  assign n213_o = {n200_o, n201_o, n202_o, n203_o};
  assign n214_o = {n204_o, n205_o, n206_o, n207_o};
  assign n215_o = {n208_o, n209_o, n210_o, n211_o};
  assign n216_o = {n212_o, n213_o, n214_o, n215_o};
  assign n217_o = data_read[31:16];
  /* TG68KdotC_Kernel.vhd:499:41  */
  assign n218_o = n195_o ? n216_o : n217_o;
  /* TG68KdotC_Kernel.vhd:497:41  */
  assign n219_o = n191_o ? last_opc_read : n218_o;
  assign n220_o = data_read[15:0];
  assign n221_o = {n219_o, n220_o};
  /* TG68KdotC_Kernel.vhd:494:25  */
  assign n222_o = n225_o ? n221_o : last_data_read;
  /* TG68KdotC_Kernel.vhd:503:61  */
  assign n223_o = last_data_in[15:0];
  /* TG68KdotC_Kernel.vhd:503:74  */
  assign n224_o = {n223_o, data_in};
  /* TG68KdotC_Kernel.vhd:494:25  */
  assign n225_o = n186_o & clkena_in;
  /* TG68KdotC_Kernel.vhd:494:25  */
  assign n226_o = clkena_in ? n224_o : last_data_in;
  /* TG68KdotC_Kernel.vhd:492:25  */
  assign n228_o = reset ? 32'b00000000000000000000000000000000 : n222_o;
  /* TG68KdotC_Kernel.vhd:492:25  */
  assign n229_o = reset ? last_data_in : n226_o;
  /* TG68KdotC_Kernel.vhd:507:65  */
  assign n233_o = memmask[1];
  /* TG68KdotC_Kernel.vhd:507:54  */
  assign n234_o = ~n233_o;
  /* TG68KdotC_Kernel.vhd:508:64  */
  assign n235_o = memread[1];
  /* TG68KdotC_Kernel.vhd:508:53  */
  assign n236_o = ~n235_o;
  /* TG68KdotC_Kernel.vhd:514:24  */
  assign n240_o = exec[40];
  /* TG68KdotC_Kernel.vhd:514:17  */
  assign n241_o = n240_o ? reg_qb : data_write_tmp;
  /* TG68KdotC_Kernel.vhd:527:39  */
  assign n242_o = addr[0];
  /* TG68KdotC_Kernel.vhd:527:34  */
  assign n243_o = oddout == n242_o;
  /* TG68KdotC_Kernel.vhd:528:61  */
  assign n245_o = {8'bX, bf_ext_out};
  /* TG68KdotC_Kernel.vhd:528:72  */
  assign n246_o = {n245_o, data_write_muxin};
  /* TG68KdotC_Kernel.vhd:530:61  */
  assign n247_o = {bf_ext_out, data_write_muxin};
  /* TG68KdotC_Kernel.vhd:530:78  */
  assign n249_o = {n247_o, 8'bX};
  /* TG68KdotC_Kernel.vhd:527:25  */
  assign n250_o = n243_o ? n246_o : n249_o;
  /* TG68KdotC_Kernel.vhd:534:30  */
  assign n251_o = memmaskmux[1];
  /* TG68KdotC_Kernel.vhd:534:33  */
  assign n252_o = ~n251_o;
  /* TG68KdotC_Kernel.vhd:535:53  */
  assign n253_o = data_write_mux[47:32];
  /* TG68KdotC_Kernel.vhd:536:33  */
  assign n254_o = memmaskmux[3];
  /* TG68KdotC_Kernel.vhd:536:36  */
  assign n255_o = ~n254_o;
  /* TG68KdotC_Kernel.vhd:537:53  */
  assign n256_o = data_write_mux[31:16];
  /* TG68KdotC_Kernel.vhd:540:38  */
  assign n257_o = memmaskmux[5:4];
  /* TG68KdotC_Kernel.vhd:540:51  */
  assign n259_o = n257_o == 2'b10;
  /* TG68KdotC_Kernel.vhd:541:61  */
  assign n260_o = data_write_mux[7:0];
  /* TG68KdotC_Kernel.vhd:541:90  */
  assign n261_o = data_write_mux[7:0];
  /* TG68KdotC_Kernel.vhd:541:74  */
  assign n262_o = {n260_o, n261_o};
  /* TG68KdotC_Kernel.vhd:542:41  */
  assign n263_o = memmaskmux[5:4];
  /* TG68KdotC_Kernel.vhd:542:54  */
  assign n265_o = n263_o == 2'b01;
  /* TG68KdotC_Kernel.vhd:543:61  */
  assign n266_o = data_write_mux[15:8];
  /* TG68KdotC_Kernel.vhd:543:91  */
  assign n267_o = data_write_mux[15:8];
  /* TG68KdotC_Kernel.vhd:543:75  */
  assign n268_o = {n266_o, n267_o};
  /* TG68KdotC_Kernel.vhd:545:61  */
  assign n269_o = data_write_mux[15:0];
  /* TG68KdotC_Kernel.vhd:542:25  */
  assign n270_o = n265_o ? n268_o : n269_o;
  /* TG68KdotC_Kernel.vhd:540:25  */
  assign n271_o = n259_o ? n262_o : n270_o;
  /* TG68KdotC_Kernel.vhd:536:17  */
  assign n272_o = n255_o ? n256_o : n271_o;
  /* TG68KdotC_Kernel.vhd:534:17  */
  assign n273_o = n252_o ? n253_o : n272_o;
  /* TG68KdotC_Kernel.vhd:548:24  */
  assign n274_o = exec[72];
  /* TG68KdotC_Kernel.vhd:549:53  */
  assign n275_o = data_write_tmp[15:8];
  /* TG68KdotC_Kernel.vhd:549:83  */
  assign n276_o = data_write_tmp[15:8];
  /* TG68KdotC_Kernel.vhd:549:67  */
  assign n277_o = {n275_o, n276_o};
  /* TG68KdotC_Kernel.vhd:548:17  */
  assign n278_o = n274_o ? n277_o : n273_o;
  /* TG68KdotC_Kernel.vhd:563:56  */
  assign n291_o = rf_dest_addr[3];
  /* TG68KdotC_Kernel.vhd:570:40  */
  assign n299_o = exec[65];
  /* TG68KdotC_Kernel.vhd:561:21  */
  assign n302_o = wwrena & clkena_lw;
  /* TG68KdotC_Kernel.vhd:561:21  */
  assign n306_o = n299_o & clkena_lw;
  /* TG68KdotC_Kernel.vhd:583:24  */
  assign n316_o = exec[30];
  /* TG68KdotC_Kernel.vhd:585:27  */
  assign n317_o = exec[62];
  /* TG68KdotC_Kernel.vhd:585:44  */
  assign n318_o = ea_only & n317_o;
  /* TG68KdotC_Kernel.vhd:587:27  */
  assign n319_o = exec[66];
  /* TG68KdotC_Kernel.vhd:589:27  */
  assign n320_o = exec[32];
  /* TG68KdotC_Kernel.vhd:594:53  */
  assign n325_o = reg_qa[15:8];
  assign n326_o = memaddr[15:8];
  assign n327_o = memaddr_a[15:8];
  assign n328_o = usp[15:8];
  assign n329_o = movec_data[15:8];
  assign n330_o = aluout[15:8];
  /* TG68KdotC_Kernel.vhd:589:17  */
  assign n331_o = n320_o ? n329_o : n330_o;
  /* TG68KdotC_Kernel.vhd:587:17  */
  assign n332_o = n319_o ? n328_o : n331_o;
  /* TG68KdotC_Kernel.vhd:585:17  */
  assign n333_o = n318_o ? n327_o : n332_o;
  /* TG68KdotC_Kernel.vhd:583:17  */
  assign n334_o = n316_o ? n326_o : n333_o;
  /* TG68KdotC_Kernel.vhd:593:17  */
  assign n335_o = bwrena ? n325_o : n334_o;
  assign n336_o = memaddr[31:16];
  assign n337_o = memaddr_a[31:16];
  assign n338_o = usp[31:16];
  assign n339_o = movec_data[31:16];
  assign n340_o = aluout[31:16];
  /* TG68KdotC_Kernel.vhd:589:17  */
  assign n341_o = n320_o ? n339_o : n340_o;
  /* TG68KdotC_Kernel.vhd:587:17  */
  assign n342_o = n319_o ? n338_o : n341_o;
  /* TG68KdotC_Kernel.vhd:585:17  */
  assign n343_o = n318_o ? n337_o : n342_o;
  /* TG68KdotC_Kernel.vhd:583:17  */
  assign n344_o = n316_o ? n336_o : n343_o;
  assign n345_o = memaddr[7:0];
  assign n346_o = memaddr_a[7:0];
  assign n347_o = usp[7:0];
  assign n348_o = movec_data[7:0];
  assign n349_o = aluout[7:0];
  /* TG68KdotC_Kernel.vhd:589:17  */
  assign n350_o = n320_o ? n348_o : n349_o;
  /* TG68KdotC_Kernel.vhd:587:17  */
  assign n351_o = n319_o ? n347_o : n350_o;
  /* TG68KdotC_Kernel.vhd:585:17  */
  assign n352_o = n318_o ? n346_o : n351_o;
  /* TG68KdotC_Kernel.vhd:583:17  */
  assign n353_o = n316_o ? n345_o : n352_o;
  /* TG68KdotC_Kernel.vhd:596:26  */
  assign n354_o = ~lwrena;
  /* TG68KdotC_Kernel.vhd:597:54  */
  assign n355_o = reg_qa[31:16];
  /* TG68KdotC_Kernel.vhd:596:17  */
  assign n356_o = n354_o ? n355_o : n344_o;
  /* TG68KdotC_Kernel.vhd:603:24  */
  assign n357_o = exec[47];
  /* TG68KdotC_Kernel.vhd:603:44  */
  assign n358_o = exec[46];
  /* TG68KdotC_Kernel.vhd:603:37  */
  assign n359_o = n357_o | n358_o;
  /* TG68KdotC_Kernel.vhd:603:65  */
  assign n360_o = exec[41];
  /* TG68KdotC_Kernel.vhd:603:58  */
  assign n361_o = n359_o | n360_o;
  /* TG68KdotC_Kernel.vhd:608:27  */
  assign n362_o = exec[34];
  /* TG68KdotC_Kernel.vhd:611:33  */
  assign n364_o = exe_datatype == 2'b00;
  /* TG68KdotC_Kernel.vhd:614:56  */
  assign n365_o = wr_areg | movem_actiond;
  /* TG68KdotC_Kernel.vhd:614:41  */
  assign n368_o = n365_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:613:33  */
  assign n370_o = exe_datatype == 2'b01;
  assign n371_o = {n370_o, n364_o};
  /* TG68KdotC_Kernel.vhd:610:25  */
  always @*
    case (n371_o)
      2'b10: n374_o = n368_o;
      2'b01: n374_o = 1'b0;
      default: n374_o = 1'b1;
    endcase
  /* TG68KdotC_Kernel.vhd:610:25  */
  always @*
    case (n371_o)
      2'b10: n377_o = 1'b0;
      2'b01: n377_o = 1'b1;
      default: n377_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:608:17  */
  assign n380_o = n362_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:608:17  */
  assign n382_o = n362_o ? n374_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:608:17  */
  assign n384_o = n362_o ? n377_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:606:17  */
  assign n386_o = regwrena_now ? 1'b1 : n380_o;
  /* TG68KdotC_Kernel.vhd:606:17  */
  assign n388_o = regwrena_now ? 1'b0 : n382_o;
  /* TG68KdotC_Kernel.vhd:606:17  */
  assign n390_o = regwrena_now ? 1'b0 : n384_o;
  /* TG68KdotC_Kernel.vhd:603:17  */
  assign n392_o = n361_o ? 1'b1 : n386_o;
  /* TG68KdotC_Kernel.vhd:603:17  */
  assign n395_o = n361_o ? 1'b1 : n388_o;
  /* TG68KdotC_Kernel.vhd:603:17  */
  assign n398_o = n361_o ? 1'b0 : n390_o;
  /* TG68KdotC_Kernel.vhd:628:24  */
  assign n403_o = exec[69];
  /* TG68KdotC_Kernel.vhd:630:26  */
  assign n404_o = set[70];
  /* TG68KdotC_Kernel.vhd:631:46  */
  assign n405_o = brief[15:12];
  /* TG68KdotC_Kernel.vhd:632:26  */
  assign n406_o = set[29];
  /* TG68KdotC_Kernel.vhd:634:59  */
  assign n407_o = sndopc[8:6];
  /* TG68KdotC_Kernel.vhd:634:52  */
  assign n409_o = {1'b0, n407_o};
  /* TG68KdotC_Kernel.vhd:639:60  */
  assign n410_o = sndopc[14:12];
  /* TG68KdotC_Kernel.vhd:639:53  */
  assign n411_o = {dest_ldrareg, n410_o};
  /* TG68KdotC_Kernel.vhd:641:55  */
  assign n412_o = last_data_read[15:12];
  /* TG68KdotC_Kernel.vhd:643:59  */
  assign n413_o = last_data_read[2:0];
  /* TG68KdotC_Kernel.vhd:643:44  */
  assign n415_o = {1'b0, n413_o};
  /* TG68KdotC_Kernel.vhd:645:51  */
  assign n416_o = sndopc[2:0];
  /* TG68KdotC_Kernel.vhd:645:44  */
  assign n418_o = {1'b0, n416_o};
  /* TG68KdotC_Kernel.vhd:649:57  */
  assign n419_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:649:50  */
  assign n420_o = {dest_areg, n419_o};
  /* TG68KdotC_Kernel.vhd:651:34  */
  assign n421_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:651:46  */
  assign n423_o = n421_o == 3'b000;
  /* TG68KdotC_Kernel.vhd:651:53  */
  assign n424_o = n423_o | data_is_source;
  /* TG68KdotC_Kernel.vhd:652:65  */
  assign n425_o = opcode[2:0];
  /* TG68KdotC_Kernel.vhd:652:58  */
  assign n426_o = {dest_areg, n425_o};
  /* TG68KdotC_Kernel.vhd:654:59  */
  assign n427_o = opcode[2:0];
  /* TG68KdotC_Kernel.vhd:654:52  */
  assign n429_o = {1'b1, n427_o};
  /* TG68KdotC_Kernel.vhd:651:25  */
  assign n430_o = n424_o ? n426_o : n429_o;
  /* TG68KdotC_Kernel.vhd:648:17  */
  assign n431_o = dest_hbits ? n420_o : n430_o;
  /* TG68KdotC_Kernel.vhd:646:17  */
  assign n433_o = setstackaddr ? 4'b1111 : n431_o;
  /* TG68KdotC_Kernel.vhd:644:17  */
  assign n434_o = dest_2ndlbits ? n418_o : n433_o;
  /* TG68KdotC_Kernel.vhd:642:17  */
  assign n435_o = dest_ldrlbits ? n415_o : n434_o;
  /* TG68KdotC_Kernel.vhd:640:17  */
  assign n436_o = dest_ldrhbits ? n412_o : n435_o;
  /* TG68KdotC_Kernel.vhd:638:17  */
  assign n437_o = dest_2ndhbits ? n411_o : n436_o;
  /* TG68KdotC_Kernel.vhd:632:17  */
  assign n438_o = n406_o ? n409_o : n437_o;
  /* TG68KdotC_Kernel.vhd:630:17  */
  assign n439_o = n404_o ? n405_o : n438_o;
  /* TG68KdotC_Kernel.vhd:628:17  */
  assign n440_o = n403_o ? rf_source_addrd : n439_o;
  /* TG68KdotC_Kernel.vhd:664:24  */
  assign n444_o = exec[69];
  /* TG68KdotC_Kernel.vhd:664:49  */
  assign n445_o = set[69];
  /* TG68KdotC_Kernel.vhd:664:43  */
  assign n446_o = n444_o | n445_o;
  /* TG68KdotC_Kernel.vhd:666:65  */
  assign n448_o = movem_regaddr ^ 4'b1111;
  /* TG68KdotC_Kernel.vhd:665:25  */
  assign n449_o = movem_presub ? n448_o : movem_regaddr;
  /* TG68KdotC_Kernel.vhd:671:53  */
  assign n450_o = sndopc[2:0];
  /* TG68KdotC_Kernel.vhd:671:46  */
  assign n452_o = {1'b0, n450_o};
  /* TG68KdotC_Kernel.vhd:673:53  */
  assign n453_o = sndopc[14:12];
  /* TG68KdotC_Kernel.vhd:673:46  */
  assign n455_o = {1'b0, n453_o};
  /* TG68KdotC_Kernel.vhd:675:53  */
  assign n456_o = sndopc[8:6];
  /* TG68KdotC_Kernel.vhd:675:46  */
  assign n458_o = {1'b0, n456_o};
  /* TG68KdotC_Kernel.vhd:677:61  */
  assign n459_o = last_data_read[2:0];
  /* TG68KdotC_Kernel.vhd:677:46  */
  assign n461_o = {1'b0, n459_o};
  /* TG68KdotC_Kernel.vhd:679:61  */
  assign n462_o = last_data_read[8:6];
  /* TG68KdotC_Kernel.vhd:679:46  */
  assign n464_o = {1'b0, n462_o};
  /* TG68KdotC_Kernel.vhd:681:61  */
  assign n465_o = opcode[2:0];
  /* TG68KdotC_Kernel.vhd:681:54  */
  assign n466_o = {source_areg, n465_o};
  /* TG68KdotC_Kernel.vhd:682:27  */
  assign n467_o = exec[36];
  /* TG68KdotC_Kernel.vhd:685:61  */
  assign n468_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:685:54  */
  assign n469_o = {source_areg, n468_o};
  /* TG68KdotC_Kernel.vhd:682:17  */
  assign n471_o = n467_o ? 4'b1111 : n469_o;
  /* TG68KdotC_Kernel.vhd:680:17  */
  assign n472_o = source_lowbits ? n466_o : n471_o;
  /* TG68KdotC_Kernel.vhd:678:17  */
  assign n473_o = source_ldrmbits ? n464_o : n472_o;
  /* TG68KdotC_Kernel.vhd:676:17  */
  assign n474_o = source_ldrlbits ? n461_o : n473_o;
  /* TG68KdotC_Kernel.vhd:674:17  */
  assign n475_o = source_2ndmbits ? n458_o : n474_o;
  /* TG68KdotC_Kernel.vhd:672:17  */
  assign n476_o = source_2ndhbits ? n455_o : n475_o;
  /* TG68KdotC_Kernel.vhd:670:17  */
  assign n477_o = source_2ndlbits ? n452_o : n476_o;
  /* TG68KdotC_Kernel.vhd:664:17  */
  assign n478_o = n446_o ? n449_o : n477_o;
  /* TG68KdotC_Kernel.vhd:695:24  */
  assign n482_o = exec[54];
  /* TG68KdotC_Kernel.vhd:697:27  */
  assign n483_o = exec[26];
  /* TG68KdotC_Kernel.vhd:697:45  */
  assign n484_o = store_in_tmp & n483_o;
  /* TG68KdotC_Kernel.vhd:699:27  */
  assign n485_o = exec[69];
  /* TG68KdotC_Kernel.vhd:699:59  */
  assign n486_o = memmaskmux[3];
  /* TG68KdotC_Kernel.vhd:699:62  */
  assign n487_o = ~n486_o;
  /* TG68KdotC_Kernel.vhd:699:46  */
  assign n488_o = n485_o | n487_o;
  /* TG68KdotC_Kernel.vhd:699:74  */
  assign n489_o = exec[39];
  /* TG68KdotC_Kernel.vhd:699:67  */
  assign n490_o = n488_o | n489_o;
  /* TG68KdotC_Kernel.vhd:699:17  */
  assign n491_o = n490_o ? addr : reg_qa;
  /* TG68KdotC_Kernel.vhd:697:17  */
  assign n492_o = n484_o ? ea_data : n491_o;
  /* TG68KdotC_Kernel.vhd:695:17  */
  assign n494_o = n482_o ? 32'b00000000000000000000000000000000 : n492_o;
  /* TG68KdotC_Kernel.vhd:710:46  */
  assign n498_o = reg_qb[15:0];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n499_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n500_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n501_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n502_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n503_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n504_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n505_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n506_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n507_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n508_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n509_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n510_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n511_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n512_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n513_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:711:58  */
  assign n514_o = op2out[15];
  assign n515_o = {n499_o, n500_o, n501_o, n502_o};
  assign n516_o = {n503_o, n504_o, n505_o, n506_o};
  assign n517_o = {n507_o, n508_o, n509_o, n510_o};
  assign n518_o = {n511_o, n512_o, n513_o, n514_o};
  assign n519_o = {n515_o, n516_o, n517_o, n518_o};
  /* TG68KdotC_Kernel.vhd:712:24  */
  assign n520_o = exec[53];
  /* TG68KdotC_Kernel.vhd:714:51  */
  assign n522_o = exec[61];
  /* TG68KdotC_Kernel.vhd:714:61  */
  assign n523_o = execopc & n522_o;
  /* TG68KdotC_Kernel.vhd:714:43  */
  assign n524_o = use_direct_data | n523_o;
  /* TG68KdotC_Kernel.vhd:714:85  */
  assign n525_o = exec[29];
  /* TG68KdotC_Kernel.vhd:714:78  */
  assign n526_o = n524_o | n525_o;
  /* TG68KdotC_Kernel.vhd:716:28  */
  assign n527_o = exec[26];
  /* TG68KdotC_Kernel.vhd:716:41  */
  assign n528_o = ~n527_o;
  /* TG68KdotC_Kernel.vhd:716:46  */
  assign n529_o = store_in_tmp & n528_o;
  /* TG68KdotC_Kernel.vhd:716:75  */
  assign n530_o = exec[27];
  /* TG68KdotC_Kernel.vhd:716:68  */
  assign n531_o = n529_o | n530_o;
  /* TG68KdotC_Kernel.vhd:718:27  */
  assign n532_o = exec[1];
  /* TG68KdotC_Kernel.vhd:719:57  */
  assign n533_o = exe_opcode[7:0];
  /* TG68KdotC_Kernel.vhd:720:69  */
  assign n534_o = exe_opcode[7];
  /* TG68KdotC_Kernel.vhd:720:69  */
  assign n535_o = exe_opcode[7];
  /* TG68KdotC_Kernel.vhd:720:69  */
  assign n536_o = exe_opcode[7];
  /* TG68KdotC_Kernel.vhd:720:69  */
  assign n537_o = exe_opcode[7];
  /* TG68KdotC_Kernel.vhd:720:69  */
  assign n538_o = exe_opcode[7];
  /* TG68KdotC_Kernel.vhd:720:69  */
  assign n539_o = exe_opcode[7];
  /* TG68KdotC_Kernel.vhd:720:69  */
  assign n540_o = exe_opcode[7];
  /* TG68KdotC_Kernel.vhd:720:69  */
  assign n541_o = exe_opcode[7];
  assign n542_o = {n534_o, n535_o, n536_o, n537_o};
  assign n543_o = {n538_o, n539_o, n540_o, n541_o};
  assign n544_o = {n542_o, n543_o};
  /* TG68KdotC_Kernel.vhd:721:27  */
  assign n545_o = exec[4];
  /* TG68KdotC_Kernel.vhd:722:57  */
  assign n546_o = exe_opcode[11:9];
  /* TG68KdotC_Kernel.vhd:723:38  */
  assign n547_o = exe_opcode[11:9];
  /* TG68KdotC_Kernel.vhd:723:51  */
  assign n549_o = n547_o == 3'b000;
  /* TG68KdotC_Kernel.vhd:723:25  */
  assign n552_o = n549_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:729:35  */
  assign n555_o = exe_datatype == 2'b10;
  /* TG68KdotC_Kernel.vhd:729:49  */
  assign n556_o = exec[11];
  /* TG68KdotC_Kernel.vhd:729:57  */
  assign n557_o = ~n556_o;
  /* TG68KdotC_Kernel.vhd:729:41  */
  assign n558_o = n557_o & n555_o;
  /* TG68KdotC_Kernel.vhd:730:55  */
  assign n559_o = reg_qb[31:16];
  /* TG68KdotC_Kernel.vhd:729:17  */
  assign n560_o = n558_o ? n559_o : n519_o;
  assign n561_o = {12'b000000000000, n552_o, n546_o};
  /* TG68KdotC_Kernel.vhd:721:17  */
  assign n562_o = n545_o ? n561_o : n498_o;
  /* TG68KdotC_Kernel.vhd:721:17  */
  assign n563_o = n545_o ? n519_o : n560_o;
  assign n564_o = {n563_o, n562_o};
  assign n565_o = {n544_o, n533_o};
  assign n566_o = n564_o[15:0];
  /* TG68KdotC_Kernel.vhd:718:17  */
  assign n567_o = n532_o ? n565_o : n566_o;
  assign n568_o = n564_o[31:16];
  /* TG68KdotC_Kernel.vhd:718:17  */
  assign n569_o = n532_o ? n519_o : n568_o;
  assign n570_o = {n569_o, n567_o};
  /* TG68KdotC_Kernel.vhd:716:17  */
  assign n571_o = n531_o ? ea_data : n570_o;
  /* TG68KdotC_Kernel.vhd:714:17  */
  assign n572_o = n526_o ? data_write_tmp : n571_o;
  assign n575_o = n572_o[31:16];
  /* TG68KdotC_Kernel.vhd:712:17  */
  assign n576_o = n520_o ? n519_o : n575_o;
  /* TG68KdotC_Kernel.vhd:732:24  */
  assign n577_o = exec[88];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n578_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n579_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n580_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n581_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n582_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n583_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n584_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n585_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n586_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n587_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n588_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n589_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n590_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n591_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n592_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n593_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n594_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n595_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n596_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n597_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n598_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n599_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n600_o = op2out[7];
  /* TG68KdotC_Kernel.vhd:733:65  */
  assign n601_o = op2out[7];
  assign n602_o = {n578_o, n579_o, n580_o, n581_o};
  assign n603_o = {n582_o, n583_o, n584_o, n585_o};
  assign n604_o = {n586_o, n587_o, n588_o, n589_o};
  assign n605_o = {n590_o, n591_o, n592_o, n593_o};
  assign n606_o = {n594_o, n595_o, n596_o, n597_o};
  assign n607_o = {n598_o, n599_o, n600_o, n601_o};
  assign n608_o = {n602_o, n603_o, n604_o, n605_o};
  assign n609_o = {n606_o, n607_o};
  assign n610_o = {n608_o, n609_o};
  assign n611_o = n521_o[15:8];
  assign n612_o = data_write_tmp[15:8];
  assign n613_o = ea_data[15:8];
  assign n614_o = n570_o[15:8];
  /* TG68KdotC_Kernel.vhd:716:17  */
  assign n615_o = n531_o ? n613_o : n614_o;
  /* TG68KdotC_Kernel.vhd:714:17  */
  assign n616_o = n526_o ? n612_o : n615_o;
  /* TG68KdotC_Kernel.vhd:712:17  */
  assign n617_o = n520_o ? n611_o : n616_o;
  assign n618_o = {n576_o, n617_o};
  /* TG68KdotC_Kernel.vhd:732:17  */
  assign n619_o = n577_o ? n610_o : n618_o;
  assign n620_o = n521_o[7:0];
  assign n621_o = data_write_tmp[7:0];
  assign n622_o = ea_data[7:0];
  assign n623_o = n570_o[7:0];
  /* TG68KdotC_Kernel.vhd:716:17  */
  assign n624_o = n531_o ? n622_o : n623_o;
  /* TG68KdotC_Kernel.vhd:714:17  */
  assign n625_o = n526_o ? n621_o : n624_o;
  /* TG68KdotC_Kernel.vhd:712:17  */
  assign n626_o = n520_o ? n620_o : n625_o;
  /* TG68KdotC_Kernel.vhd:753:40  */
  assign n631_o = exec[82];
  /* TG68KdotC_Kernel.vhd:753:33  */
  assign n633_o = n631_o ? 1'b1 : use_direct_data;
  /* TG68KdotC_Kernel.vhd:759:56  */
  assign n634_o = set[27];
  /* TG68KdotC_Kernel.vhd:759:50  */
  assign n635_o = endopc | n634_o;
  /* TG68KdotC_Kernel.vhd:759:33  */
  assign n637_o = n635_o ? 1'b0 : n633_o;
  /* TG68KdotC_Kernel.vhd:756:33  */
  assign n639_o = set_direct_data ? 1'b1 : n637_o;
  /* TG68KdotC_Kernel.vhd:756:33  */
  assign n642_o = set_direct_data ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:762:56  */
  assign n644_o = set_exec[0];
  /* TG68KdotC_Kernel.vhd:769:41  */
  assign n646_o = set_z_error ? 1'b1 : z_error;
  /* TG68KdotC_Kernel.vhd:772:52  */
  assign n647_o = set_exec[0];
  /* TG68KdotC_Kernel.vhd:772:75  */
  assign n649_o = state == 2'b11;
  /* TG68KdotC_Kernel.vhd:772:66  */
  assign n650_o = n649_o & n647_o;
  /* TG68KdotC_Kernel.vhd:772:41  */
  assign n652_o = n650_o ? 1'b1 : n639_o;
  /* TG68KdotC_Kernel.vhd:776:49  */
  assign n654_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:776:62  */
  assign n655_o = exec[80];
  /* TG68KdotC_Kernel.vhd:776:55  */
  assign n656_o = n654_o | n655_o;
  /* TG68KdotC_Kernel.vhd:776:41  */
  assign n658_o = n656_o ? 1'b1 : store_in_tmp;
  /* TG68KdotC_Kernel.vhd:779:69  */
  assign n660_o = state == 2'b00;
  /* TG68KdotC_Kernel.vhd:779:60  */
  assign n661_o = n660_o & direct_data;
  /* TG68KdotC_Kernel.vhd:779:41  */
  assign n663_o = n661_o ? 1'b1 : n658_o;
  /* TG68KdotC_Kernel.vhd:764:33  */
  assign n665_o = endopc ? 1'b0 : n663_o;
  /* TG68KdotC_Kernel.vhd:764:33  */
  assign n667_o = endopc ? 1'b0 : writepcnext;
  /* TG68KdotC_Kernel.vhd:764:33  */
  assign n668_o = endopc ? n639_o : n652_o;
  /* TG68KdotC_Kernel.vhd:764:33  */
  assign n670_o = endopc ? 1'b0 : n646_o;
  /* TG68KdotC_Kernel.vhd:784:41  */
  assign n672_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:784:55  */
  assign n673_o = exec[79];
  /* TG68KdotC_Kernel.vhd:784:69  */
  assign n674_o = ~n673_o;
  /* TG68KdotC_Kernel.vhd:784:47  */
  assign n675_o = n674_o & n672_o;
  /* TG68KdotC_Kernel.vhd:786:43  */
  assign n676_o = exec[71];
  /* TG68KdotC_Kernel.vhd:788:43  */
  assign n677_o = exec[44];
  /* TG68KdotC_Kernel.vhd:788:92  */
  assign n679_o = state == 2'b00;
  /* TG68KdotC_Kernel.vhd:788:83  */
  assign n680_o = n679_o & direct_data;
  /* TG68KdotC_Kernel.vhd:788:63  */
  assign n681_o = n677_o | n680_o;
  /* TG68KdotC_Kernel.vhd:788:33  */
  assign n682_o = n681_o ? last_data_read : ea_data;
  /* TG68KdotC_Kernel.vhd:786:33  */
  assign n683_o = n676_o ? addr : n682_o;
  /* TG68KdotC_Kernel.vhd:784:33  */
  assign n684_o = n675_o ? data_read : n683_o;
  /* TG68KdotC_Kernel.vhd:794:43  */
  assign n685_o = exec[25];
  /* TG68KdotC_Kernel.vhd:797:50  */
  assign n687_o = $unsigned(micro_state) >= $unsigned(7'b0110111);
  /* TG68KdotC_Kernel.vhd:797:74  */
  assign n689_o = $unsigned(micro_state) <= $unsigned(7'b0111101);
  /* TG68KdotC_Kernel.vhd:797:58  */
  assign n690_o = n689_o & n687_o;
  /* TG68KdotC_Kernel.vhd:799:50  */
  assign n692_o = micro_state == 7'b0110010;
  /* TG68KdotC_Kernel.vhd:802:66  */
  assign n693_o = trap_trap | trap_trapv;
  /* TG68KdotC_Kernel.vhd:802:87  */
  assign n694_o = exec[43];
  /* TG68KdotC_Kernel.vhd:802:80  */
  assign n695_o = n693_o | n694_o;
  /* TG68KdotC_Kernel.vhd:802:98  */
  assign n696_o = n695_o | z_error;
  /* TG68KdotC_Kernel.vhd:803:51  */
  assign n698_o = micro_state == 7'b0110011;
  /* TG68KdotC_Kernel.vhd:809:100  */
  assign n699_o = trap_vector[11:0];
  /* TG68KdotC_Kernel.vhd:809:87  */
  assign n701_o = {4'b0010, n699_o};
  /* TG68KdotC_Kernel.vhd:811:61  */
  assign n702_o = trap_berr | trap_addr_error;
  /* TG68KdotC_Kernel.vhd:812:100  */
  assign n703_o = trap_vector[11:0];
  /* TG68KdotC_Kernel.vhd:812:87  */
  assign n705_o = {4'b1111, n703_o};
  /* TG68KdotC_Kernel.vhd:813:74  */
  assign n706_o = trap_trap | trap_trapv;
  /* TG68KdotC_Kernel.vhd:813:95  */
  assign n707_o = exec[43];
  /* TG68KdotC_Kernel.vhd:813:88  */
  assign n708_o = n706_o | n707_o;
  /* TG68KdotC_Kernel.vhd:813:106  */
  assign n709_o = n708_o | z_error;
  /* TG68KdotC_Kernel.vhd:815:100  */
  assign n710_o = trap_vector[11:0];
  /* TG68KdotC_Kernel.vhd:815:87  */
  assign n712_o = {4'b0000, n710_o};
  /* TG68KdotC_Kernel.vhd:816:74  */
  assign n713_o = trap_trap | trap_trapv;
  /* TG68KdotC_Kernel.vhd:816:95  */
  assign n714_o = exec[43];
  /* TG68KdotC_Kernel.vhd:816:88  */
  assign n715_o = n713_o | n714_o;
  /* TG68KdotC_Kernel.vhd:816:106  */
  assign n716_o = n715_o | z_error;
  /* TG68KdotC_Kernel.vhd:811:41  */
  assign n717_o = n702_o ? n705_o : n712_o;
  /* TG68KdotC_Kernel.vhd:811:41  */
  assign n718_o = n702_o ? n709_o : n716_o;
  /* TG68KdotC_Kernel.vhd:807:41  */
  assign n719_o = usestackframe2 ? n701_o : n717_o;
  /* TG68KdotC_Kernel.vhd:807:41  */
  assign n720_o = usestackframe2 ? n667_o : n718_o;
  /* TG68KdotC_Kernel.vhd:821:43  */
  assign n721_o = exec[64];
  /* TG68KdotC_Kernel.vhd:823:43  */
  assign n722_o = exec[61];
  /* TG68KdotC_Kernel.vhd:825:43  */
  assign n723_o = exec[62];
  /* TG68KdotC_Kernel.vhd:825:60  */
  assign n724_o = ea_only & n723_o;
  /* TG68KdotC_Kernel.vhd:829:65  */
  assign n726_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:829:56  */
  assign n727_o = n726_o & exec_direct;
  /* TG68KdotC_Kernel.vhd:831:49  */
  assign n728_o = exec[37];
  /* TG68KdotC_Kernel.vhd:832:94  */
  assign n729_o = data_write_tmp[23:0];
  assign n730_o = data_read[31:8];
  /* TG68KdotC_Kernel.vhd:831:41  */
  assign n731_o = n728_o ? n729_o : n730_o;
  assign n732_o = data_read[7:0];
  /* TG68KdotC_Kernel.vhd:834:43  */
  assign n733_o = exec[37];
  /* TG68KdotC_Kernel.vhd:835:78  */
  assign n734_o = reg_qb[31:16];
  /* TG68KdotC_Kernel.vhd:839:91  */
  assign n735_o = {trap_sr, flags};
  assign n736_o = op2out[15:0];
  /* TG68KdotC_Kernel.vhd:838:33  */
  assign n737_o = writesr ? n735_o : n736_o;
  assign n738_o = op2out[31:16];
  assign n739_o = data_write_tmp[31:16];
  /* TG68KdotC_Kernel.vhd:838:33  */
  assign n740_o = writesr ? n739_o : n738_o;
  assign n741_o = {n740_o, n737_o};
  /* TG68KdotC_Kernel.vhd:836:33  */
  assign n742_o = direct_data ? last_data_read : n741_o;
  assign n743_o = n742_o[15:0];
  /* TG68KdotC_Kernel.vhd:834:33  */
  assign n744_o = n733_o ? n734_o : n743_o;
  assign n745_o = n742_o[31:16];
  assign n746_o = data_write_tmp[31:16];
  /* TG68KdotC_Kernel.vhd:834:33  */
  assign n747_o = n733_o ? n746_o : n745_o;
  assign n748_o = {n747_o, n744_o};
  assign n749_o = {n731_o, n732_o};
  /* TG68KdotC_Kernel.vhd:829:33  */
  assign n750_o = n727_o ? n749_o : n748_o;
  /* TG68KdotC_Kernel.vhd:827:33  */
  assign n751_o = execopc ? aluout : n750_o;
  /* TG68KdotC_Kernel.vhd:825:33  */
  assign n752_o = n724_o ? addr : n751_o;
  /* TG68KdotC_Kernel.vhd:823:33  */
  assign n753_o = n722_o ? op1out : n752_o;
  /* TG68KdotC_Kernel.vhd:821:33  */
  assign n754_o = n721_o ? data_write_tmp : n753_o;
  assign n755_o = n754_o[15:0];
  /* TG68KdotC_Kernel.vhd:803:33  */
  assign n756_o = n698_o ? n719_o : n755_o;
  assign n757_o = n754_o[31:16];
  assign n758_o = data_write_tmp[31:16];
  /* TG68KdotC_Kernel.vhd:803:33  */
  assign n759_o = n698_o ? n758_o : n757_o;
  /* TG68KdotC_Kernel.vhd:803:33  */
  assign n760_o = n698_o ? n720_o : n667_o;
  assign n761_o = {n759_o, n756_o};
  /* TG68KdotC_Kernel.vhd:799:33  */
  assign n762_o = n692_o ? exe_pc : n761_o;
  /* TG68KdotC_Kernel.vhd:799:33  */
  assign n763_o = n692_o ? n696_o : n760_o;
  /* TG68KdotC_Kernel.vhd:799:33  */
  assign n766_o = n692_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:797:33  */
  assign n768_o = n690_o ? 32'b00000000000000000000000000000000 : n762_o;
  /* TG68KdotC_Kernel.vhd:797:33  */
  assign n769_o = n690_o ? n667_o : n763_o;
  /* TG68KdotC_Kernel.vhd:797:33  */
  assign n771_o = n690_o ? 1'b0 : n766_o;
  /* TG68KdotC_Kernel.vhd:794:33  */
  assign n772_o = n685_o ? tg68_pc_add : n768_o;
  /* TG68KdotC_Kernel.vhd:794:33  */
  assign n773_o = n685_o ? n667_o : n769_o;
  /* TG68KdotC_Kernel.vhd:794:33  */
  assign n775_o = n685_o ? 1'b0 : n771_o;
  /* TG68KdotC_Kernel.vhd:792:33  */
  assign n776_o = writepc ? tg68_pc : n772_o;
  /* TG68KdotC_Kernel.vhd:792:33  */
  assign n777_o = writepc ? n667_o : n773_o;
  /* TG68KdotC_Kernel.vhd:792:33  */
  assign n779_o = writepc ? 1'b0 : n775_o;
  /* TG68KdotC_Kernel.vhd:750:25  */
  assign n781_o = clkena_lw ? n684_o : ea_data;
  /* TG68KdotC_Kernel.vhd:750:25  */
  assign n782_o = clkena_lw ? n776_o : data_write_tmp;
  /* TG68KdotC_Kernel.vhd:750:25  */
  assign n783_o = clkena_lw ? n665_o : store_in_tmp;
  /* TG68KdotC_Kernel.vhd:750:25  */
  assign n784_o = clkena_lw ? n777_o : writepcnext;
  /* TG68KdotC_Kernel.vhd:750:25  */
  assign n785_o = clkena_lw ? n644_o : exec_direct;
  /* TG68KdotC_Kernel.vhd:750:25  */
  assign n786_o = clkena_lw ? n668_o : use_direct_data;
  /* TG68KdotC_Kernel.vhd:750:25  */
  assign n787_o = clkena_lw ? n642_o : direct_data;
  /* TG68KdotC_Kernel.vhd:750:25  */
  assign n788_o = clkena_lw ? n779_o : usestackframe2;
  /* TG68KdotC_Kernel.vhd:750:25  */
  assign n789_o = clkena_lw ? n670_o : z_error;
  /* TG68KdotC_Kernel.vhd:744:25  */
  assign n790_o = reset ? ea_data : n781_o;
  /* TG68KdotC_Kernel.vhd:744:25  */
  assign n791_o = reset ? data_write_tmp : n782_o;
  /* TG68KdotC_Kernel.vhd:744:25  */
  assign n793_o = reset ? 1'b0 : n783_o;
  /* TG68KdotC_Kernel.vhd:744:25  */
  assign n795_o = reset ? 1'b0 : n784_o;
  /* TG68KdotC_Kernel.vhd:744:25  */
  assign n796_o = reset ? exec_direct : n785_o;
  /* TG68KdotC_Kernel.vhd:744:25  */
  assign n798_o = reset ? 1'b0 : n786_o;
  /* TG68KdotC_Kernel.vhd:744:25  */
  assign n800_o = reset ? 1'b0 : n787_o;
  /* TG68KdotC_Kernel.vhd:744:25  */
  assign n801_o = reset ? usestackframe2 : n788_o;
  /* TG68KdotC_Kernel.vhd:744:25  */
  assign n803_o = reset ? 1'b0 : n789_o;
  /* TG68KdotC_Kernel.vhd:852:25  */
  assign n816_o = brief[11];
  /* TG68KdotC_Kernel.vhd:853:46  */
  assign n817_o = op1out[31:16];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n818_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n819_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n820_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n821_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n822_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n823_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n824_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n825_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n826_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n827_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n828_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n829_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n830_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n831_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n832_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:855:55  */
  assign n833_o = op1out[15];
  assign n834_o = {n818_o, n819_o, n820_o, n821_o};
  assign n835_o = {n822_o, n823_o, n824_o, n825_o};
  assign n836_o = {n826_o, n827_o, n828_o, n829_o};
  assign n837_o = {n830_o, n831_o, n832_o, n833_o};
  assign n838_o = {n834_o, n835_o, n836_o, n837_o};
  /* TG68KdotC_Kernel.vhd:852:17  */
  assign n839_o = n816_o ? n817_o : n838_o;
  /* TG68KdotC_Kernel.vhd:857:48  */
  assign n840_o = op1out[15:0];
  /* TG68KdotC_Kernel.vhd:857:41  */
  assign n841_o = {op1outbrief, n840_o};
  /* TG68KdotC_Kernel.vhd:858:42  */
  assign n842_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:858:50  */
  assign n844_o = 1'b1 & n842_o;
  /* TG68KdotC_Kernel.vhd:858:35  */
  assign n846_o = 1'b0 | n844_o;
  /* TG68KdotC_Kernel.vhd:859:35  */
  assign n847_o = brief[10:9];
  /* TG68KdotC_Kernel.vhd:860:77  */
  assign n848_o = op1out[15:0];
  /* TG68KdotC_Kernel.vhd:860:70  */
  assign n849_o = {op1outbrief, n848_o};
  /* TG68KdotC_Kernel.vhd:860:33  */
  assign n851_o = n847_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:861:70  */
  assign n852_o = op1outbrief[14:0];
  /* TG68KdotC_Kernel.vhd:861:90  */
  assign n853_o = op1out[15:0];
  /* TG68KdotC_Kernel.vhd:861:83  */
  assign n854_o = {n852_o, n853_o};
  /* TG68KdotC_Kernel.vhd:861:103  */
  assign n856_o = {n854_o, 1'b0};
  /* TG68KdotC_Kernel.vhd:861:33  */
  assign n858_o = n847_o == 2'b01;
  /* TG68KdotC_Kernel.vhd:862:70  */
  assign n859_o = op1outbrief[13:0];
  /* TG68KdotC_Kernel.vhd:862:90  */
  assign n860_o = op1out[15:0];
  /* TG68KdotC_Kernel.vhd:862:83  */
  assign n861_o = {n859_o, n860_o};
  /* TG68KdotC_Kernel.vhd:862:103  */
  assign n863_o = {n861_o, 2'b00};
  /* TG68KdotC_Kernel.vhd:862:33  */
  assign n865_o = n847_o == 2'b10;
  /* TG68KdotC_Kernel.vhd:863:70  */
  assign n866_o = op1outbrief[12:0];
  /* TG68KdotC_Kernel.vhd:863:90  */
  assign n867_o = op1out[15:0];
  /* TG68KdotC_Kernel.vhd:863:83  */
  assign n868_o = {n866_o, n867_o};
  /* TG68KdotC_Kernel.vhd:863:103  */
  assign n870_o = {n868_o, 3'b000};
  /* TG68KdotC_Kernel.vhd:863:33  */
  assign n872_o = n847_o == 2'b11;
  assign n873_o = {n872_o, n865_o, n858_o, n851_o};
  /* TG68KdotC_Kernel.vhd:859:25  */
  always @*
    case (n873_o)
      4'b1000: n874_o = n870_o;
      4'b0100: n874_o = n863_o;
      4'b0010: n874_o = n856_o;
      4'b0001: n874_o = n849_o;
      default: n874_o = n841_o;
    endcase
  /* TG68KdotC_Kernel.vhd:858:17  */
  assign n875_o = n846_o ? n874_o : n841_o;
  assign n882_o = trap_vector[9:0];
  /* TG68KdotC_Kernel.vhd:879:33  */
  assign n883_o = trap_berr ? 10'b0000001000 : n882_o;
  /* TG68KdotC_Kernel.vhd:882:33  */
  assign n885_o = trap_addr_error ? 10'b0000001100 : n883_o;
  /* TG68KdotC_Kernel.vhd:885:33  */
  assign n887_o = trap_illegal ? 10'b0000010000 : n885_o;
  /* TG68KdotC_Kernel.vhd:888:33  */
  assign n889_o = set_z_error ? 10'b0000010100 : n887_o;
  /* TG68KdotC_Kernel.vhd:891:40  */
  assign n890_o = exec[43];
  /* TG68KdotC_Kernel.vhd:891:33  */
  assign n892_o = n890_o ? 10'b0000011000 : n889_o;
  /* TG68KdotC_Kernel.vhd:894:33  */
  assign n894_o = trap_trapv ? 10'b0000011100 : n892_o;
  /* TG68KdotC_Kernel.vhd:897:33  */
  assign n896_o = trap_priv ? 10'b0000100000 : n894_o;
  /* TG68KdotC_Kernel.vhd:900:33  */
  assign n898_o = trap_trace ? 10'b0000100100 : n896_o;
  /* TG68KdotC_Kernel.vhd:903:33  */
  assign n900_o = trap_1010 ? 10'b0000101000 : n898_o;
  /* TG68KdotC_Kernel.vhd:906:33  */
  assign n902_o = trap_1111 ? 10'b0000101100 : n900_o;
  /* TG68KdotC_Kernel.vhd:910:83  */
  assign n903_o = opcode[3:0];
  /* TG68KdotC_Kernel.vhd:910:75  */
  assign n905_o = {4'b0010, n903_o};
  /* TG68KdotC_Kernel.vhd:910:96  */
  assign n907_o = {n905_o, 2'b00};
  /* TG68KdotC_Kernel.vhd:909:33  */
  assign n908_o = trap_trap ? n907_o : n902_o;
  /* TG68KdotC_Kernel.vhd:912:55  */
  assign n909_o = trap_interrupt | set_vectoraddr;
  /* TG68KdotC_Kernel.vhd:913:76  */
  assign n911_o = {ipl_vec, 2'b00};
  /* TG68KdotC_Kernel.vhd:912:33  */
  assign n912_o = n909_o ? n911_o : n908_o;
  assign n913_o = {22'b0000000000000000000000, n912_o};
  /* TG68KdotC_Kernel.vhd:918:55  */
  assign n916_o = trap_vector + vbr;
  /* TG68KdotC_Kernel.vhd:917:17  */
  assign n917_o = use_vbr_stackframe ? n916_o : trap_vector;
  /* TG68KdotC_Kernel.vhd:924:60  */
  assign n919_o = memaddr_a[4];
  /* TG68KdotC_Kernel.vhd:924:60  */
  assign n920_o = memaddr_a[4];
  /* TG68KdotC_Kernel.vhd:924:60  */
  assign n921_o = memaddr_a[4];
  assign n922_o = {n919_o, n920_o, n921_o};
  /* TG68KdotC_Kernel.vhd:925:61  */
  assign n923_o = memaddr_a[7];
  /* TG68KdotC_Kernel.vhd:925:61  */
  assign n924_o = memaddr_a[7];
  /* TG68KdotC_Kernel.vhd:925:61  */
  assign n925_o = memaddr_a[7];
  /* TG68KdotC_Kernel.vhd:925:61  */
  assign n926_o = memaddr_a[7];
  /* TG68KdotC_Kernel.vhd:925:61  */
  assign n927_o = memaddr_a[7];
  /* TG68KdotC_Kernel.vhd:925:61  */
  assign n928_o = memaddr_a[7];
  /* TG68KdotC_Kernel.vhd:925:61  */
  assign n929_o = memaddr_a[7];
  /* TG68KdotC_Kernel.vhd:925:61  */
  assign n930_o = memaddr_a[7];
  assign n931_o = {n923_o, n924_o, n925_o, n926_o};
  assign n932_o = {n927_o, n928_o, n929_o, n930_o};
  assign n933_o = {n931_o, n932_o};
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n934_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n935_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n936_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n937_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n938_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n939_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n940_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n941_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n942_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n943_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n944_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n945_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n946_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n947_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n948_o = memaddr_a[15];
  /* TG68KdotC_Kernel.vhd:926:62  */
  assign n949_o = memaddr_a[15];
  assign n950_o = {n934_o, n935_o, n936_o, n937_o};
  assign n951_o = {n938_o, n939_o, n940_o, n941_o};
  assign n952_o = {n942_o, n943_o, n944_o, n945_o};
  assign n953_o = {n946_o, n947_o, n948_o, n949_o};
  assign n954_o = {n950_o, n951_o, n952_o, n953_o};
  /* TG68KdotC_Kernel.vhd:928:32  */
  assign n955_o = exec[70];
  /* TG68KdotC_Kernel.vhd:929:55  */
  assign n956_o = briefdata + memaddr_delta;
  /* TG68KdotC_Kernel.vhd:931:72  */
  assign n957_o = last_data_read[7:0];
  assign n958_o = last_data_read[7:0];
  /* TG68KdotC_Kernel.vhd:930:25  */
  assign n959_o = setdispbyte ? n957_o : n958_o;
  assign n960_o = last_data_read[31:8];
  assign n961_o = {n954_o, n933_o};
  /* TG68KdotC_Kernel.vhd:930:25  */
  assign n962_o = setdispbyte ? n961_o : n960_o;
  assign n963_o = {n962_o, n959_o};
  /* TG68KdotC_Kernel.vhd:928:25  */
  assign n964_o = n955_o ? n956_o : n963_o;
  /* TG68KdotC_Kernel.vhd:935:26  */
  assign n965_o = set[47];
  /* TG68KdotC_Kernel.vhd:936:31  */
  assign n966_o = set[73];
  /* TG68KdotC_Kernel.vhd:938:39  */
  assign n969_o = datatype == 2'b00;
  /* TG68KdotC_Kernel.vhd:938:52  */
  assign n970_o = set[50];
  /* TG68KdotC_Kernel.vhd:938:60  */
  assign n971_o = ~n970_o;
  /* TG68KdotC_Kernel.vhd:938:45  */
  assign n972_o = n971_o & n969_o;
  /* TG68KdotC_Kernel.vhd:938:25  */
  assign n975_o = n972_o ? 5'b11111 : 5'b11110;
  /* TG68KdotC_Kernel.vhd:936:25  */
  assign n976_o = n966_o ? 5'b11100 : n975_o;
  /* TG68KdotC_Kernel.vhd:944:53  */
  assign n978_o = {1'b1, ripl_nr};
  /* TG68KdotC_Kernel.vhd:944:61  */
  assign n980_o = {n978_o, 1'b0};
  /* TG68KdotC_Kernel.vhd:943:17  */
  assign n981_o = interrupt ? n980_o : 5'b00000;
  /* TG68KdotC_Kernel.vhd:935:17  */
  assign n982_o = n965_o ? n976_o : n981_o;
  assign n983_o = n964_o[4:0];
  /* TG68KdotC_Kernel.vhd:927:17  */
  assign n984_o = setdisp ? n983_o : n982_o;
  assign n985_o = n964_o[31:5];
  assign n986_o = {n954_o, n933_o, n922_o};
  /* TG68KdotC_Kernel.vhd:927:17  */
  assign n987_o = setdisp ? n985_o : n986_o;
  /* TG68KdotC_Kernel.vhd:949:40  */
  assign n989_o = exec[71];
  /* TG68KdotC_Kernel.vhd:949:66  */
  assign n991_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:949:83  */
  assign n992_o = memread[0];
  /* TG68KdotC_Kernel.vhd:949:72  */
  assign n993_o = n992_o & n991_o;
  /* TG68KdotC_Kernel.vhd:949:57  */
  assign n994_o = n989_o | n993_o;
  /* TG68KdotC_Kernel.vhd:954:46  */
  assign n996_o = memmaskmux[3];
  /* TG68KdotC_Kernel.vhd:954:49  */
  assign n997_o = ~n996_o;
  /* TG68KdotC_Kernel.vhd:954:61  */
  assign n998_o = exec[55];
  /* TG68KdotC_Kernel.vhd:954:54  */
  assign n999_o = n997_o | n998_o;
  /* TG68KdotC_Kernel.vhd:956:42  */
  assign n1000_o = set[83];
  /* TG68KdotC_Kernel.vhd:958:43  */
  assign n1001_o = exec[58];
  /* TG68KdotC_Kernel.vhd:960:43  */
  assign n1002_o = exec[63];
  /* TG68KdotC_Kernel.vhd:960:70  */
  assign n1004_o = setstate == 2'b00;
  /* TG68KdotC_Kernel.vhd:960:58  */
  assign n1005_o = n1004_o & n1002_o;
  /* TG68KdotC_Kernel.vhd:962:42  */
  assign n1006_o = set[45];
  /* TG68KdotC_Kernel.vhd:964:47  */
  assign n1008_o = setstate == 2'b00;
  /* TG68KdotC_Kernel.vhd:966:43  */
  assign n1009_o = exec[22];
  /* TG68KdotC_Kernel.vhd:973:53  */
  assign n1010_o = ~interrupt;
  /* TG68KdotC_Kernel.vhd:973:75  */
  assign n1011_o = ~suppress_base;
  /* TG68KdotC_Kernel.vhd:973:58  */
  assign n1012_o = n1011_o & n1010_o;
  /* TG68KdotC_Kernel.vhd:973:41  */
  assign n1015_o = n1012_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:969:33  */
  assign n1016_o = set_vectoraddr ? trap_vector_vbr : memaddr_a;
  /* TG68KdotC_Kernel.vhd:969:33  */
  assign n1018_o = set_vectoraddr ? 1'b0 : n1015_o;
  /* TG68KdotC_Kernel.vhd:966:33  */
  assign n1019_o = n1009_o ? ea_data : n1016_o;
  /* TG68KdotC_Kernel.vhd:966:33  */
  assign n1021_o = n1009_o ? memaddr_a : 32'b00000000000000000000000000000000;
  /* TG68KdotC_Kernel.vhd:966:33  */
  assign n1023_o = n1009_o ? 1'b0 : n1018_o;
  /* TG68KdotC_Kernel.vhd:964:33  */
  assign n1024_o = n1008_o ? tg68_pc_add : n1019_o;
  /* TG68KdotC_Kernel.vhd:964:33  */
  assign n1026_o = n1008_o ? 32'b00000000000000000000000000000000 : n1021_o;
  /* TG68KdotC_Kernel.vhd:964:33  */
  assign n1028_o = n1008_o ? 1'b0 : n1023_o;
  /* TG68KdotC_Kernel.vhd:962:33  */
  assign n1029_o = n1006_o ? last_data_read : n1024_o;
  /* TG68KdotC_Kernel.vhd:962:33  */
  assign n1031_o = n1006_o ? 32'b00000000000000000000000000000000 : n1026_o;
  /* TG68KdotC_Kernel.vhd:962:33  */
  assign n1033_o = n1006_o ? 1'b0 : n1028_o;
  /* TG68KdotC_Kernel.vhd:960:33  */
  assign n1034_o = n1005_o ? addr : n1029_o;
  /* TG68KdotC_Kernel.vhd:960:33  */
  assign n1036_o = n1005_o ? 32'b00000000000000000000000000000000 : n1031_o;
  /* TG68KdotC_Kernel.vhd:960:33  */
  assign n1038_o = n1005_o ? 1'b0 : n1033_o;
  /* TG68KdotC_Kernel.vhd:958:33  */
  assign n1039_o = n1001_o ? data_read : n1034_o;
  /* TG68KdotC_Kernel.vhd:958:33  */
  assign n1041_o = n1001_o ? 32'b00000000000000000000000000000000 : n1036_o;
  /* TG68KdotC_Kernel.vhd:958:33  */
  assign n1043_o = n1001_o ? 1'b0 : n1038_o;
  /* TG68KdotC_Kernel.vhd:956:33  */
  assign n1044_o = n1000_o ? tmp_tg68_pc : n1039_o;
  /* TG68KdotC_Kernel.vhd:956:33  */
  assign n1046_o = n1000_o ? 32'b00000000000000000000000000000000 : n1041_o;
  /* TG68KdotC_Kernel.vhd:956:33  */
  assign n1048_o = n1000_o ? 1'b0 : n1043_o;
  /* TG68KdotC_Kernel.vhd:954:33  */
  assign n1049_o = n999_o ? addsub_q : n1044_o;
  /* TG68KdotC_Kernel.vhd:954:33  */
  assign n1051_o = n999_o ? 32'b00000000000000000000000000000000 : n1046_o;
  /* TG68KdotC_Kernel.vhd:954:33  */
  assign n1054_o = n999_o ? 1'b0 : n1048_o;
  /* TG68KdotC_Kernel.vhd:981:53  */
  assign n1056_o = memread[0];
  /* TG68KdotC_Kernel.vhd:981:73  */
  assign n1057_o = state[1];
  /* TG68KdotC_Kernel.vhd:981:64  */
  assign n1058_o = n1057_o & n1056_o;
  /* TG68KdotC_Kernel.vhd:981:100  */
  assign n1059_o = ~movem_presub;
  /* TG68KdotC_Kernel.vhd:981:84  */
  assign n1060_o = n1058_o | n1059_o;
  /* TG68KdotC_Kernel.vhd:948:25  */
  assign n1062_o = n994_o & clkena_in;
  /* TG68KdotC_Kernel.vhd:948:25  */
  assign n1063_o = n1060_o & clkena_in;
  /* TG68KdotC_Kernel.vhd:987:53  */
  assign n1072_o = memaddr_delta_rega + memaddr_delta_regb;
  /* TG68KdotC_Kernel.vhd:989:36  */
  assign n1073_o = memaddr_reg + memaddr_delta;
  /* TG68KdotC_Kernel.vhd:990:41  */
  assign n1074_o = memaddr_reg + memaddr_delta;
  /* TG68KdotC_Kernel.vhd:992:28  */
  assign n1075_o = ~use_base;
  /* TG68KdotC_Kernel.vhd:992:17  */
  assign n1077_o = n1075_o ? 32'b00000000000000000000000000000000 : reg_qa;
  /* TG68KdotC_Kernel.vhd:1007:17  */
  assign n1081_o = tg68_pc_brw ? tmp_tg68_pc : tg68_pc;
  /* TG68KdotC_Kernel.vhd:1012:40  */
  assign n1083_o = pc_datab[2];
  /* TG68KdotC_Kernel.vhd:1013:60  */
  assign n1084_o = pc_datab[3];
  /* TG68KdotC_Kernel.vhd:1013:60  */
  assign n1085_o = pc_datab[3];
  /* TG68KdotC_Kernel.vhd:1013:60  */
  assign n1086_o = pc_datab[3];
  /* TG68KdotC_Kernel.vhd:1013:60  */
  assign n1087_o = pc_datab[3];
  assign n1088_o = {n1084_o, n1085_o, n1086_o, n1087_o};
  /* TG68KdotC_Kernel.vhd:1014:61  */
  assign n1089_o = pc_datab[7];
  /* TG68KdotC_Kernel.vhd:1014:61  */
  assign n1090_o = pc_datab[7];
  /* TG68KdotC_Kernel.vhd:1014:61  */
  assign n1091_o = pc_datab[7];
  /* TG68KdotC_Kernel.vhd:1014:61  */
  assign n1092_o = pc_datab[7];
  /* TG68KdotC_Kernel.vhd:1014:61  */
  assign n1093_o = pc_datab[7];
  /* TG68KdotC_Kernel.vhd:1014:61  */
  assign n1094_o = pc_datab[7];
  /* TG68KdotC_Kernel.vhd:1014:61  */
  assign n1095_o = pc_datab[7];
  /* TG68KdotC_Kernel.vhd:1014:61  */
  assign n1096_o = pc_datab[7];
  assign n1097_o = {n1089_o, n1090_o, n1091_o, n1092_o};
  assign n1098_o = {n1093_o, n1094_o, n1095_o, n1096_o};
  assign n1099_o = {n1097_o, n1098_o};
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1100_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1101_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1102_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1103_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1104_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1105_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1106_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1107_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1108_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1109_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1110_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1111_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1112_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1113_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1114_o = pc_datab[15];
  /* TG68KdotC_Kernel.vhd:1015:62  */
  assign n1115_o = pc_datab[15];
  assign n1116_o = {n1100_o, n1101_o, n1102_o, n1103_o};
  assign n1117_o = {n1104_o, n1105_o, n1106_o, n1107_o};
  assign n1118_o = {n1108_o, n1109_o, n1110_o, n1111_o};
  assign n1119_o = {n1112_o, n1113_o, n1114_o, n1115_o};
  assign n1120_o = {n1116_o, n1117_o, n1118_o, n1119_o};
  assign n1124_o = n1082_o[0];
  /* TG68KdotC_Kernel.vhd:1019:24  */
  assign n1125_o = exec[25];
  assign n1129_o = n1121_o[0];
  assign n1130_o = n1082_o[1];
  /* TG68KdotC_Kernel.vhd:1016:17  */
  assign n1131_o = interrupt ? n1129_o : n1130_o;
  /* TG68KdotC_Kernel.vhd:1020:25  */
  assign n1132_o = writepcbig ? 1'b1 : n1131_o;
  assign n1133_o = n1121_o[1];
  assign n1134_o = n1082_o[2];
  /* TG68KdotC_Kernel.vhd:1016:17  */
  assign n1135_o = interrupt ? n1133_o : n1134_o;
  /* TG68KdotC_Kernel.vhd:1020:25  */
  assign n1136_o = writepcbig ? n1135_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1020:25  */
  assign n1137_o = writepcbig ? 1'b1 : n1083_o;
  /* TG68KdotC_Kernel.vhd:1026:47  */
  assign n1138_o = ~use_vbr_stackframe;
  /* TG68KdotC_Kernel.vhd:1026:71  */
  assign n1139_o = trap_trap | trap_trapv;
  /* TG68KdotC_Kernel.vhd:1026:96  */
  assign n1140_o = exec[43];
  /* TG68KdotC_Kernel.vhd:1026:89  */
  assign n1141_o = n1139_o | n1140_o;
  /* TG68KdotC_Kernel.vhd:1026:111  */
  assign n1142_o = n1141_o | z_error;
  /* TG68KdotC_Kernel.vhd:1026:52  */
  assign n1143_o = n1142_o & n1138_o;
  /* TG68KdotC_Kernel.vhd:1026:128  */
  assign n1144_o = n1143_o | writepcnext;
  /* TG68KdotC_Kernel.vhd:1026:25  */
  assign n1146_o = n1144_o ? 1'b1 : n1132_o;
  /* TG68KdotC_Kernel.vhd:1029:28  */
  assign n1148_o = state == 2'b00;
  assign n1150_o = n1121_o[0];
  assign n1151_o = n1082_o[1];
  /* TG68KdotC_Kernel.vhd:1016:17  */
  assign n1152_o = interrupt ? n1150_o : n1151_o;
  /* TG68KdotC_Kernel.vhd:1029:17  */
  assign n1153_o = n1148_o ? 1'b1 : n1152_o;
  assign n1154_o = {n1137_o, n1136_o, n1146_o};
  assign n1155_o = n1154_o[0];
  /* TG68KdotC_Kernel.vhd:1019:17  */
  assign n1156_o = n1125_o ? n1155_o : n1153_o;
  assign n1157_o = n1154_o[2:1];
  assign n1158_o = n1121_o[1];
  assign n1159_o = n1082_o[2];
  /* TG68KdotC_Kernel.vhd:1016:17  */
  assign n1160_o = interrupt ? n1158_o : n1159_o;
  assign n1161_o = {n1083_o, n1160_o};
  /* TG68KdotC_Kernel.vhd:1019:17  */
  assign n1162_o = n1125_o ? n1157_o : n1161_o;
  /* TG68KdotC_Kernel.vhd:1036:63  */
  assign n1166_o = opcode[7:0];
  assign n1167_o = last_data_read[7:0];
  /* TG68KdotC_Kernel.vhd:1033:25  */
  assign n1168_o = tg68_pc_word ? n1167_o : n1166_o;
  assign n1169_o = last_data_read[31:8];
  assign n1170_o = {n1120_o, n1099_o};
  /* TG68KdotC_Kernel.vhd:1033:25  */
  assign n1171_o = tg68_pc_word ? n1169_o : n1170_o;
  assign n1172_o = {n1171_o, n1168_o};
  assign n1173_o = {n1120_o, n1099_o, n1088_o, n1162_o, n1156_o, n1124_o};
  /* TG68KdotC_Kernel.vhd:1032:17  */
  assign n1174_o = tg68_pc_brw ? n1172_o : n1173_o;
  /* TG68KdotC_Kernel.vhd:1040:40  */
  assign n1175_o = pc_dataa + pc_datab;
  /* TG68KdotC_Kernel.vhd:1045:28  */
  assign n1177_o = setstate == 2'b00;
  /* TG68KdotC_Kernel.vhd:1045:54  */
  assign n1179_o = next_micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:1045:34  */
  assign n1180_o = n1179_o & n1177_o;
  /* TG68KdotC_Kernel.vhd:1045:75  */
  assign n1181_o = ~setnextpass;
  /* TG68KdotC_Kernel.vhd:1045:60  */
  assign n1182_o = n1181_o & n1180_o;
  /* TG68KdotC_Kernel.vhd:1045:100  */
  assign n1183_o = ~exec_write_back;
  /* TG68KdotC_Kernel.vhd:1045:113  */
  assign n1185_o = state == 2'b11;
  /* TG68KdotC_Kernel.vhd:1045:105  */
  assign n1186_o = n1183_o | n1185_o;
  /* TG68KdotC_Kernel.vhd:1045:80  */
  assign n1187_o = n1186_o & n1182_o;
  /* TG68KdotC_Kernel.vhd:1045:135  */
  assign n1189_o = set_rot_cnt == 6'b000001;
  /* TG68KdotC_Kernel.vhd:1045:120  */
  assign n1190_o = n1189_o & n1187_o;
  /* TG68KdotC_Kernel.vhd:1045:157  */
  assign n1191_o = set_exec[31];
  /* TG68KdotC_Kernel.vhd:1045:165  */
  assign n1192_o = ~n1191_o;
  /* TG68KdotC_Kernel.vhd:1045:145  */
  assign n1193_o = n1192_o & n1190_o;
  /* TG68KdotC_Kernel.vhd:1047:35  */
  assign n1194_o = flagssr[2:0];
  /* TG68KdotC_Kernel.vhd:1047:47  */
  assign n1195_o = $unsigned(n1194_o) < $unsigned(ipl_nr);
  /* TG68KdotC_Kernel.vhd:1047:64  */
  assign n1197_o = ipl_nr == 3'b111;
  /* TG68KdotC_Kernel.vhd:1047:55  */
  assign n1198_o = n1195_o | n1197_o;
  /* TG68KdotC_Kernel.vhd:1047:72  */
  assign n1199_o = n1198_o | make_trace;
  /* TG68KdotC_Kernel.vhd:1047:90  */
  assign n1200_o = n1199_o | make_berr;
  /* TG68KdotC_Kernel.vhd:1049:35  */
  assign n1201_o = ~stop;
  /* TG68KdotC_Kernel.vhd:1049:25  */
  assign n1204_o = n1201_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1047:25  */
  assign n1206_o = n1200_o ? 1'b0 : n1204_o;
  /* TG68KdotC_Kernel.vhd:1047:25  */
  assign n1209_o = n1200_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1045:17  */
  assign n1211_o = n1193_o ? n1206_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1045:17  */
  assign n1215_o = n1193_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1045:17  */
  assign n1218_o = n1193_o ? n1209_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1054:28  */
  assign n1221_o = setstate == 2'b00;
  /* TG68KdotC_Kernel.vhd:1054:54  */
  assign n1223_o = next_micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:1054:34  */
  assign n1224_o = n1223_o & n1221_o;
  /* TG68KdotC_Kernel.vhd:1054:79  */
  assign n1225_o = ~set_direct_data;
  /* TG68KdotC_Kernel.vhd:1054:60  */
  assign n1226_o = n1225_o & n1224_o;
  /* TG68KdotC_Kernel.vhd:1054:104  */
  assign n1227_o = ~exec_write_back;
  /* TG68KdotC_Kernel.vhd:1054:118  */
  assign n1229_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:1054:137  */
  assign n1230_o = ~addrvalue;
  /* TG68KdotC_Kernel.vhd:1054:124  */
  assign n1231_o = n1230_o & n1229_o;
  /* TG68KdotC_Kernel.vhd:1054:109  */
  assign n1232_o = n1227_o | n1231_o;
  /* TG68KdotC_Kernel.vhd:1054:84  */
  assign n1233_o = n1232_o & n1226_o;
  /* TG68KdotC_Kernel.vhd:1054:17  */
  assign n1236_o = n1233_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1058:27  */
  assign n1238_o = ~ipl;
  /* TG68KdotC_Kernel.vhd:1088:59  */
  assign n1240_o = memmask[3:0];
  /* TG68KdotC_Kernel.vhd:1088:71  */
  assign n1242_o = {n1240_o, 2'b11};
  /* TG68KdotC_Kernel.vhd:1089:59  */
  assign n1243_o = memread[1:0];
  /* TG68KdotC_Kernel.vhd:1089:82  */
  assign n1244_o = memmaskmux[5:4];
  /* TG68KdotC_Kernel.vhd:1089:71  */
  assign n1245_o = {n1243_o, n1244_o};
  /* TG68KdotC_Kernel.vhd:1093:48  */
  assign n1246_o = exec[57];
  /* TG68KdotC_Kernel.vhd:1095:51  */
  assign n1247_o = exec[63];
  /* TG68KdotC_Kernel.vhd:1097:54  */
  assign n1249_o = state == 2'b00;
  /* TG68KdotC_Kernel.vhd:1097:60  */
  assign n1250_o = n1249_o | tg68_pc_brw;
  /* TG68KdotC_Kernel.vhd:1097:90  */
  assign n1251_o = ~stop;
  /* TG68KdotC_Kernel.vhd:1097:82  */
  assign n1252_o = n1251_o & n1250_o;
  /* TG68KdotC_Kernel.vhd:1097:41  */
  assign n1253_o = n1252_o ? tg68_pc_add : tg68_pc;
  /* TG68KdotC_Kernel.vhd:1095:41  */
  assign n1254_o = n1247_o ? addr : n1253_o;
  /* TG68KdotC_Kernel.vhd:1093:41  */
  assign n1255_o = n1246_o ? data_read : n1254_o;
  /* TG68KdotC_Kernel.vhd:1087:33  */
  assign n1256_o = clkena_in ? n1255_o : tg68_pc;
  /* TG68KdotC_Kernel.vhd:1087:33  */
  assign n1257_o = clkena_in ? n1242_o : memmask;
  /* TG68KdotC_Kernel.vhd:1087:33  */
  assign n1258_o = clkena_in ? n1245_o : memread;
  /* TG68KdotC_Kernel.vhd:1115:53  */
  assign n1259_o = ~trap_berr;
  /* TG68KdotC_Kernel.vhd:1116:68  */
  assign n1260_o = berr | make_berr;
  /* TG68KdotC_Kernel.vhd:1115:41  */
  assign n1262_o = n1259_o ? n1260_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1121:71  */
  assign n1263_o = ~setinterrupt;
  /* TG68KdotC_Kernel.vhd:1121:67  */
  assign n1264_o = n1263_o & stop;
  /* TG68KdotC_Kernel.vhd:1121:58  */
  assign n1265_o = set_stop | n1264_o;
  /* TG68KdotC_Kernel.vhd:1134:75  */
  assign n1267_o = {5'b00011, ipl_nr};
  /* TG68KdotC_Kernel.vhd:1130:49  */
  assign n1270_o = make_berr ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1130:49  */
  assign n1273_o = make_berr ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1130:49  */
  assign n1274_o = make_berr ? ripl_nr : ipl_nr;
  /* TG68KdotC_Kernel.vhd:1130:49  */
  assign n1275_o = make_berr ? ipl_vec : n1267_o;
  /* TG68KdotC_Kernel.vhd:1128:49  */
  assign n1277_o = make_trace ? 1'b0 : n1270_o;
  /* TG68KdotC_Kernel.vhd:1128:49  */
  assign n1281_o = make_trace ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1128:49  */
  assign n1284_o = make_trace ? 1'b0 : n1273_o;
  /* TG68KdotC_Kernel.vhd:1128:49  */
  assign n1286_o = make_trace ? ripl_nr : n1274_o;
  /* TG68KdotC_Kernel.vhd:1128:49  */
  assign n1287_o = make_trace ? ipl_vec : n1275_o;
  /* TG68KdotC_Kernel.vhd:1122:41  */
  assign n1288_o = setinterrupt ? n1277_o : trap_berr;
  /* TG68KdotC_Kernel.vhd:1122:41  */
  assign n1289_o = setinterrupt ? n1281_o : trap_trace;
  /* TG68KdotC_Kernel.vhd:1122:41  */
  assign n1290_o = setinterrupt ? n1284_o : trap_interrupt;
  /* TG68KdotC_Kernel.vhd:1122:41  */
  assign n1292_o = setinterrupt ? 1'b0 : n1262_o;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1293_o = n1496_o ? n1286_o : ripl_nr;
  /* TG68KdotC_Kernel.vhd:1122:41  */
  assign n1294_o = setinterrupt ? n1287_o : ipl_vec;
  /* TG68KdotC_Kernel.vhd:1138:55  */
  assign n1296_o = micro_state == 7'b0110011;
  /* TG68KdotC_Kernel.vhd:1138:80  */
  assign n1297_o = ~ipl_autovector;
  /* TG68KdotC_Kernel.vhd:1138:62  */
  assign n1298_o = n1297_o & n1296_o;
  /* TG68KdotC_Kernel.vhd:1139:74  */
  assign n1299_o = last_data_read[7:0];
  /* TG68KdotC_Kernel.vhd:1138:41  */
  assign n1300_o = n1298_o ? n1299_o : n1294_o;
  /* TG68KdotC_Kernel.vhd:1141:49  */
  assign n1302_o = state == 2'b00;
  /* TG68KdotC_Kernel.vhd:1142:75  */
  assign n1303_o = data_read[15:0];
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1304_o = n1478_o ? tg68_pc : last_opc_pc;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1305_o = n1479_o ? n1303_o : last_opc_read;
  /* TG68KdotC_Kernel.vhd:1150:53  */
  assign n1306_o = opcode[7:0];
  /* TG68KdotC_Kernel.vhd:1150:65  */
  assign n1308_o = n1306_o == 8'b00000000;
  /* TG68KdotC_Kernel.vhd:1150:86  */
  assign n1309_o = opcode[7:0];
  /* TG68KdotC_Kernel.vhd:1150:98  */
  assign n1311_o = n1309_o == 8'b11111111;
  /* TG68KdotC_Kernel.vhd:1150:77  */
  assign n1312_o = n1308_o | n1311_o;
  /* TG68KdotC_Kernel.vhd:1150:110  */
  assign n1313_o = n1312_o | data_is_source;
  /* TG68KdotC_Kernel.vhd:1150:41  */
  assign n1315_o = n1313_o ? 1'b1 : tg68_pc_word;
  /* TG68KdotC_Kernel.vhd:1145:41  */
  assign n1317_o = setopcode ? 1'b0 : n1315_o;
  /* TG68KdotC_Kernel.vhd:1145:41  */
  assign n1319_o = setopcode ? 1'b0 : n1288_o;
  /* TG68KdotC_Kernel.vhd:1145:41  */
  assign n1321_o = setopcode ? 1'b0 : n1289_o;
  /* TG68KdotC_Kernel.vhd:1145:41  */
  assign n1323_o = setopcode ? 1'b0 : n1290_o;
  /* TG68KdotC_Kernel.vhd:1154:48  */
  assign n1324_o = exec[29];
  /* TG68KdotC_Kernel.vhd:1158:84  */
  assign n1325_o = {26'b0, bf_width};  //  uext
  /* TG68KdotC_Kernel.vhd:1158:84  */
  assign n1326_o = bf_full_offset + n1325_o;
  /* TG68KdotC_Kernel.vhd:1158:93  */
  assign n1328_o = n1326_o + 32'b00000000000000000000000000000001;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1329_o = n1505_o ? bf_width : alu_width;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1330_o = n1506_o ? bf_shift : alu_bf_shift;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1331_o = n1507_o ? n1328_o : alu_bf_ffo_offset;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1332_o = n1508_o ? bf_loffset : alu_bf_loffset;
  /* TG68KdotC_Kernel.vhd:1161:62  */
  assign n1333_o = setstate[1];
  /* TG68KdotC_Kernel.vhd:1161:50  */
  assign n1334_o = ~n1333_o;
  /* TG68KdotC_Kernel.vhd:1161:93  */
  assign n1335_o = setstate[0];
  /* TG68KdotC_Kernel.vhd:1161:81  */
  assign n1336_o = ~n1335_o;
  /* TG68KdotC_Kernel.vhd:1161:77  */
  assign n1337_o = pcbase & n1336_o;
  /* TG68KdotC_Kernel.vhd:1161:66  */
  assign n1338_o = n1334_o | n1337_o;
  /* TG68KdotC_Kernel.vhd:1162:58  */
  assign n1339_o = setstate[1];
  /* TG68KdotC_Kernel.vhd:1162:67  */
  assign n1340_o = ~pcbase;
  /* TG68KdotC_Kernel.vhd:1162:89  */
  assign n1341_o = setstate[0];
  /* TG68KdotC_Kernel.vhd:1162:78  */
  assign n1342_o = n1340_o | n1341_o;
  /* TG68KdotC_Kernel.vhd:1162:62  */
  assign n1343_o = n1339_o & n1342_o;
  assign n1345_o = {n1338_o, n1343_o};
  /* TG68KdotC_Kernel.vhd:1163:41  */
  assign n1346_o = interrupt ? 2'b11 : n1345_o;
  /* TG68KdotC_Kernel.vhd:1167:49  */
  assign n1348_o = state == 2'b11;
  /* TG68KdotC_Kernel.vhd:1169:55  */
  assign n1350_o = setstate == 2'b10;
  /* TG68KdotC_Kernel.vhd:1169:77  */
  assign n1351_o = ~setaddrvalue;
  /* TG68KdotC_Kernel.vhd:1169:61  */
  assign n1352_o = n1351_o & n1350_o;
  /* TG68KdotC_Kernel.vhd:1169:82  */
  assign n1353_o = write_back & n1352_o;
  /* TG68KdotC_Kernel.vhd:1169:41  */
  assign n1355_o = n1353_o ? 1'b1 : exec_write_back;
  /* TG68KdotC_Kernel.vhd:1167:41  */
  assign n1357_o = n1348_o ? 1'b0 : n1355_o;
  /* TG68KdotC_Kernel.vhd:1172:50  */
  assign n1359_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:1172:69  */
  assign n1360_o = ~addrvalue;
  /* TG68KdotC_Kernel.vhd:1172:56  */
  assign n1361_o = n1360_o & n1359_o;
  /* TG68KdotC_Kernel.vhd:1172:74  */
  assign n1362_o = write_back & n1361_o;
  /* TG68KdotC_Kernel.vhd:1172:105  */
  assign n1364_o = setstate != 2'b10;
  /* TG68KdotC_Kernel.vhd:1172:93  */
  assign n1365_o = n1364_o & n1362_o;
  /* TG68KdotC_Kernel.vhd:1172:127  */
  assign n1367_o = set_rot_cnt != 6'b000001;
  /* TG68KdotC_Kernel.vhd:1172:113  */
  assign n1368_o = n1365_o | n1367_o;
  /* TG68KdotC_Kernel.vhd:1172:164  */
  assign n1369_o = ~interrupt;
  /* TG68KdotC_Kernel.vhd:1172:151  */
  assign n1370_o = n1369_o & stop;
  /* TG68KdotC_Kernel.vhd:1172:138  */
  assign n1371_o = n1368_o | n1370_o;
  /* TG68KdotC_Kernel.vhd:1172:181  */
  assign n1372_o = set_exec[31];
  /* TG68KdotC_Kernel.vhd:1172:170  */
  assign n1373_o = n1371_o | n1372_o;
  /* TG68KdotC_Kernel.vhd:1176:59  */
  assign n1374_o = exec_write_back & execopc;
  /* TG68KdotC_Kernel.vhd:1184:60  */
  assign n1377_o = setstate == 2'b01;
  /* TG68KdotC_Kernel.vhd:1187:59  */
  assign n1378_o = exec[29];
  /* TG68KdotC_Kernel.vhd:1191:58  */
  assign n1379_o = set[73];
  /* TG68KdotC_Kernel.vhd:1196:67  */
  assign n1381_o = set_datatype == 2'b00;
  /* TG68KdotC_Kernel.vhd:1196:85  */
  assign n1382_o = setstate[1];
  /* TG68KdotC_Kernel.vhd:1196:73  */
  assign n1383_o = n1382_o & n1381_o;
  /* TG68KdotC_Kernel.vhd:1199:63  */
  assign n1384_o = set[72];
  /* TG68KdotC_Kernel.vhd:1199:57  */
  assign n1387_o = n1384_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1196:49  */
  assign n1390_o = n1383_o ? 6'b101111 : 6'b100111;
  /* TG68KdotC_Kernel.vhd:1196:49  */
  assign n1393_o = n1383_o ? 6'b101111 : 6'b100111;
  /* TG68KdotC_Kernel.vhd:1196:49  */
  assign n1395_o = n1383_o ? n1387_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1191:49  */
  assign n1397_o = n1379_o ? 6'b100001 : n1390_o;
  /* TG68KdotC_Kernel.vhd:1191:49  */
  assign n1399_o = n1379_o ? 6'b100001 : n1393_o;
  /* TG68KdotC_Kernel.vhd:1191:49  */
  assign n1401_o = n1379_o ? 1'b0 : n1395_o;
  /* TG68KdotC_Kernel.vhd:1187:49  */
  assign n1402_o = n1378_o ? set_memmask : n1397_o;
  /* TG68KdotC_Kernel.vhd:1187:49  */
  assign n1403_o = n1378_o ? set_memmask : n1399_o;
  /* TG68KdotC_Kernel.vhd:1187:49  */
  assign n1404_o = n1378_o ? set_oddout : n1401_o;
  /* TG68KdotC_Kernel.vhd:1184:49  */
  assign n1406_o = n1377_o ? 6'b111111 : n1402_o;
  /* TG68KdotC_Kernel.vhd:1184:49  */
  assign n1408_o = n1377_o ? 6'b111111 : n1403_o;
  /* TG68KdotC_Kernel.vhd:1184:49  */
  assign n1409_o = n1377_o ? oddout : n1404_o;
  /* TG68KdotC_Kernel.vhd:1176:41  */
  assign n1410_o = n1374_o ? 2'b01 : n1346_o;
  /* TG68KdotC_Kernel.vhd:1176:41  */
  assign n1412_o = n1374_o ? 2'b11 : setstate;
  /* TG68KdotC_Kernel.vhd:1176:41  */
  assign n1414_o = n1374_o ? 1'b0 : setaddrvalue;
  /* TG68KdotC_Kernel.vhd:1176:41  */
  assign n1415_o = n1374_o ? wbmemmask : n1406_o;
  /* TG68KdotC_Kernel.vhd:1176:41  */
  assign n1416_o = n1374_o ? wbmemmask : n1408_o;
  /* TG68KdotC_Kernel.vhd:1176:41  */
  assign n1417_o = n1374_o ? oddout : n1409_o;
  /* TG68KdotC_Kernel.vhd:1172:41  */
  assign n1418_o = n1373_o ? n1346_o : n1410_o;
  /* TG68KdotC_Kernel.vhd:1172:41  */
  assign n1420_o = n1373_o ? 2'b01 : n1412_o;
  /* TG68KdotC_Kernel.vhd:1172:41  */
  assign n1422_o = n1373_o ? 1'b0 : n1414_o;
  /* TG68KdotC_Kernel.vhd:1172:41  */
  assign n1424_o = n1373_o ? 6'b111111 : n1415_o;
  /* TG68KdotC_Kernel.vhd:1172:41  */
  assign n1425_o = n1373_o ? wbmemmask : n1416_o;
  /* TG68KdotC_Kernel.vhd:1172:41  */
  assign n1426_o = n1373_o ? oddout : n1417_o;
  /* TG68KdotC_Kernel.vhd:1215:78  */
  assign n1427_o = set_writepcbig | writepcbig;
  /* TG68KdotC_Kernel.vhd:1211:41  */
  assign n1429_o = decodeopc ? 1'b0 : n1427_o;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1430_o = n1488_o ? set_rot_bits : rot_bits;
  /* TG68KdotC_Kernel.vhd:1217:65  */
  assign n1431_o = exec[24];
  /* TG68KdotC_Kernel.vhd:1217:58  */
  assign n1432_o = decodeopc | n1431_o;
  /* TG68KdotC_Kernel.vhd:1217:92  */
  assign n1434_o = rot_cnt != 6'b000001;
  /* TG68KdotC_Kernel.vhd:1217:82  */
  assign n1435_o = n1432_o | n1434_o;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1436_o = n1489_o ? set_rot_cnt : rot_cnt;
  /* TG68KdotC_Kernel.vhd:1223:55  */
  assign n1437_o = setstate[1];
  /* TG68KdotC_Kernel.vhd:1223:86  */
  assign n1438_o = set[62];
  /* TG68KdotC_Kernel.vhd:1223:79  */
  assign n1439_o = n1438_o & ea_only;
  /* TG68KdotC_Kernel.vhd:1223:63  */
  assign n1440_o = n1437_o | n1439_o;
  /* TG68KdotC_Kernel.vhd:1223:41  */
  assign n1442_o = n1440_o ? 1'b0 : suppress_base;
  /* TG68KdotC_Kernel.vhd:1221:41  */
  assign n1444_o = set_suppress_base ? 1'b1 : n1442_o;
  /* TG68KdotC_Kernel.vhd:1227:57  */
  assign n1445_o = state[1];
  /* TG68KdotC_Kernel.vhd:1230:75  */
  assign n1446_o = data_read[15:0];
  /* TG68KdotC_Kernel.vhd:1227:49  */
  assign n1447_o = n1445_o ? last_opc_read : n1446_o;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1448_o = n1482_o ? n1447_o : brief;
  /* TG68KdotC_Kernel.vhd:1234:66  */
  assign n1449_o = ~berr;
  /* TG68KdotC_Kernel.vhd:1234:58  */
  assign n1450_o = n1449_o & setopcode;
  /* TG68KdotC_Kernel.vhd:1235:57  */
  assign n1452_o = state == 2'b00;
  /* TG68KdotC_Kernel.vhd:1236:76  */
  assign n1453_o = data_read[15:0];
  /* TG68KdotC_Kernel.vhd:1235:49  */
  assign n1454_o = n1452_o ? n1453_o : last_opc_read;
  /* TG68KdotC_Kernel.vhd:1235:49  */
  assign n1455_o = n1452_o ? tg68_pc : last_opc_pc;
  /* TG68KdotC_Kernel.vhd:1243:64  */
  assign n1456_o = setinterrupt | setopcode;
  /* TG68KdotC_Kernel.vhd:1248:68  */
  assign n1457_o = setnextpass | regdirectsource;
  /* TG68KdotC_Kernel.vhd:1248:49  */
  assign n1459_o = n1457_o ? 1'b1 : nextpass;
  /* TG68KdotC_Kernel.vhd:1243:41  */
  assign n1461_o = n1456_o ? 16'b0100111001110001 : opcode;
  /* TG68KdotC_Kernel.vhd:1243:41  */
  assign n1463_o = n1456_o ? 1'b0 : n1459_o;
  /* TG68KdotC_Kernel.vhd:1234:41  */
  assign n1464_o = n1450_o ? n1454_o : n1461_o;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1465_o = n1477_o ? n1455_o : exe_pc;
  /* TG68KdotC_Kernel.vhd:1234:41  */
  assign n1467_o = n1450_o ? 1'b0 : n1463_o;
  /* TG68KdotC_Kernel.vhd:1253:58  */
  assign n1468_o = decodeopc | interrupt;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1469_o = n1493_o ? flagssr : trap_sr;
  assign n1470_o = n9781_o[1:0];
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1471_o = clkena_lw ? n1418_o : n1470_o;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1472_o = clkena_lw ? n1420_o : state;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1473_o = clkena_lw ? set_datatype : exe_datatype;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1474_o = clkena_lw ? n1422_o : addrvalue;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1475_o = clkena_lw ? n1464_o : opcode;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1476_o = clkena_lw ? opcode : exe_opcode;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1477_o = n1450_o & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1478_o = n1302_o & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1479_o = n1302_o & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1480_o = clkena_lw ? n1467_o : nextpass;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1481_o = clkena_lw ? n1317_o : tg68_pc_word;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1482_o = getbrief & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1483_o = clkena_lw ? n1357_o : exec_write_back;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1484_o = clkena_lw ? n1429_o : writepcbig;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1485_o = clkena_lw ? setopcode : decodeopc;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1486_o = clkena_lw ? setexecopc : execopc;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1487_o = clkena_lw ? setendopc : endopc;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1488_o = decodeopc & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1489_o = n1435_o & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1490_o = clkena_lw ? n1319_o : trap_berr;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1491_o = clkena_lw ? n1321_o : trap_trace;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1492_o = clkena_lw ? n1323_o : trap_interrupt;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1493_o = n1468_o & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1494_o = clkena_lw ? n1292_o : make_berr;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1495_o = clkena_lw ? n1265_o : stop;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1496_o = setinterrupt & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1497_o = clkena_lw ? n1300_o : ipl_vec;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1498_o = clkena_lw ? setinterrupt : interrupt;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1499_o = clkena_lw ? n1444_o : suppress_base;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1500_o = clkena_lw ? n1424_o : n1257_o;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1502_o = clkena_lw ? 4'b1111 : n1258_o;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1503_o = clkena_lw ? n1425_o : wbmemmask;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1504_o = clkena_lw ? n1426_o : oddout;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1505_o = n1324_o & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1506_o = n1324_o & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1507_o = n1324_o & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1101:33  */
  assign n1508_o = n1324_o & clkena_lw;
  assign n1509_o = n9781_o[1:0];
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1510_o = reset ? n1509_o : n1471_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1512_o = reset ? 32'b00000000000000000000000000000100 : n1256_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1514_o = reset ? 2'b01 : n1472_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1515_o = reset ? exe_datatype : n1473_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1517_o = reset ? 1'b0 : n1474_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1519_o = reset ? 16'b0010111001111001 : n1475_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1520_o = reset ? exe_opcode : n1476_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1521_o = reset ? exe_pc : n1465_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1522_o = reset ? last_opc_pc : n1304_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1524_o = reset ? 16'b0100111011111001 : n1305_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1525_o = reset ? nextpass : n1480_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1527_o = reset ? 1'b0 : n1481_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1528_o = reset ? brief : n1448_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1530_o = reset ? 1'b0 : n1483_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1532_o = reset ? 1'b0 : n1484_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1534_o = reset ? 1'b0 : n1485_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1536_o = reset ? 1'b0 : n1486_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1538_o = reset ? 1'b0 : n1487_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1539_o = reset ? rot_bits : n1430_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1541_o = reset ? 6'b000001 : n1436_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1543_o = reset ? 1'b0 : n1490_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1545_o = reset ? 1'b0 : n1491_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1547_o = reset ? 1'b0 : n1492_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1548_o = reset ? trap_sr : n1469_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1550_o = reset ? 1'b0 : n1494_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1552_o = reset ? 1'b0 : n1495_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1553_o = reset ? ripl_nr : n1293_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1554_o = reset ? ipl_vec : n1497_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1556_o = reset ? 1'b0 : n1498_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1558_o = reset ? 1'b0 : n1499_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1560_o = reset ? 6'b111111 : n1500_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1561_o = reset ? memread : n1502_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1562_o = reset ? wbmemmask : n1503_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1563_o = reset ? oddout : n1504_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1564_o = reset ? alu_width : n1329_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1565_o = reset ? alu_bf_shift : n1330_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1566_o = reset ? alu_bf_ffo_offset : n1331_o;
  /* TG68KdotC_Kernel.vhd:1060:25  */
  assign n1567_o = reset ? alu_bf_loffset : n1332_o;
  /* TG68KdotC_Kernel.vhd:1264:54  */
  assign n1608_o = set_pcbase | pcbase;
  /* TG68KdotC_Kernel.vhd:1265:60  */
  assign n1609_o = state[1];
  /* TG68KdotC_Kernel.vhd:1265:81  */
  assign n1610_o = ~movem_run;
  /* TG68KdotC_Kernel.vhd:1265:68  */
  assign n1611_o = n1610_o & n1609_o;
  /* TG68KdotC_Kernel.vhd:1265:51  */
  assign n1612_o = setexecopc | n1611_o;
  /* TG68KdotC_Kernel.vhd:1265:33  */
  assign n1614_o = n1612_o ? 1'b0 : n1608_o;
  /* TG68KdotC_Kernel.vhd:1263:25  */
  assign n1615_o = clkena_lw ? n1614_o : pcbase;
  /* TG68KdotC_Kernel.vhd:1261:25  */
  assign n1617_o = reset ? 1'b1 : n1615_o;
  /* TG68KdotC_Kernel.vhd:1271:54  */
  assign n1618_o = set[0];
  /* TG68KdotC_Kernel.vhd:1271:70  */
  assign n1619_o = set[85];
  /* TG68KdotC_Kernel.vhd:1271:64  */
  assign n1620_o = n1618_o | n1619_o;
  /* TG68KdotC_Kernel.vhd:1272:58  */
  assign n1623_o = set[3];
  /* TG68KdotC_Kernel.vhd:1272:73  */
  assign n1624_o = set[86];
  /* TG68KdotC_Kernel.vhd:1272:67  */
  assign n1625_o = n1623_o | n1624_o;
  assign n1626_o = set[88:87];
  /* TG68KdotC_Kernel.vhd:1274:52  */
  assign n1627_o = set[47];
  /* TG68KdotC_Kernel.vhd:1274:67  */
  assign n1628_o = set[48];
  /* TG68KdotC_Kernel.vhd:1274:61  */
  assign n1629_o = n1627_o | n1628_o;
  assign n1630_o = set[84:49];
  assign n1631_o = set[47:0];
  /* TG68KdotC_Kernel.vhd:1276:58  */
  assign n1632_o = set_exec | set;
  /* TG68KdotC_Kernel.vhd:1277:67  */
  assign n1633_o = set_exec[0];
  /* TG68KdotC_Kernel.vhd:1277:83  */
  assign n1634_o = set[0];
  /* TG68KdotC_Kernel.vhd:1277:77  */
  assign n1635_o = n1633_o | n1634_o;
  /* TG68KdotC_Kernel.vhd:1277:99  */
  assign n1636_o = set[85];
  /* TG68KdotC_Kernel.vhd:1277:93  */
  assign n1637_o = n1635_o | n1636_o;
  assign n1639_o = n1632_o[84:0];
  /* TG68KdotC_Kernel.vhd:1278:71  */
  assign n1640_o = set_exec[3];
  /* TG68KdotC_Kernel.vhd:1278:86  */
  assign n1641_o = set[3];
  /* TG68KdotC_Kernel.vhd:1278:80  */
  assign n1642_o = n1640_o | n1641_o;
  /* TG68KdotC_Kernel.vhd:1278:101  */
  assign n1643_o = set[86];
  /* TG68KdotC_Kernel.vhd:1278:95  */
  assign n1644_o = n1642_o | n1643_o;
  assign n1645_o = n1632_o[88:87];
  /* TG68KdotC_Kernel.vhd:1275:33  */
  assign n1647_o = setexecopc ? set_exec_tas : 1'b0;
  assign n1649_o = {n1645_o, n1644_o, n1637_o, n1639_o};
  assign n1650_o = {n1626_o, n1625_o, n1620_o, n1630_o, n1629_o, n1631_o};
  /* TG68KdotC_Kernel.vhd:1281:56  */
  assign n1652_o = set[71];
  /* TG68KdotC_Kernel.vhd:1281:69  */
  assign n1653_o = n1652_o | setopcode;
  assign n1654_o = n1649_o[88:72];
  assign n1655_o = n1650_o[88:72];
  /* TG68KdotC_Kernel.vhd:1275:33  */
  assign n1656_o = setexecopc ? n1654_o : n1655_o;
  assign n1657_o = n1649_o[70:0];
  assign n1658_o = n1650_o[70:0];
  /* TG68KdotC_Kernel.vhd:1275:33  */
  assign n1659_o = setexecopc ? n1657_o : n1658_o;
  assign n1661_o = {n1656_o, n1653_o, n1659_o};
  /* TG68KdotC_Kernel.vhd:1291:26  */
  assign n1669_o = sndopc[11];
  /* TG68KdotC_Kernel.vhd:1292:48  */
  assign n1670_o = reg_qa[4:0];
  /* TG68KdotC_Kernel.vhd:1292:41  */
  assign n1672_o = {1'b0, n1670_o};
  /* TG68KdotC_Kernel.vhd:1294:48  */
  assign n1673_o = sndopc[10:6];
  /* TG68KdotC_Kernel.vhd:1294:41  */
  assign n1675_o = {1'b0, n1673_o};
  /* TG68KdotC_Kernel.vhd:1296:26  */
  assign n1677_o = sndopc[11];
  /* TG68KdotC_Kernel.vhd:1300:61  */
  assign n1678_o = sndopc[10:6];
  assign n1680_o = n1679_o[31:5];
  assign n1681_o = {n1680_o, n1678_o};
  /* TG68KdotC_Kernel.vhd:1296:17  */
  assign n1682_o = n1677_o ? reg_qa : n1681_o;
  /* TG68KdotC_Kernel.vhd:1304:26  */
  assign n1684_o = sndopc[5];
  /* TG68KdotC_Kernel.vhd:1305:55  */
  assign n1685_o = reg_qb[4:0];
  /* TG68KdotC_Kernel.vhd:1305:67  */
  assign n1687_o = n1685_o - 5'b00001;
  /* TG68KdotC_Kernel.vhd:1307:55  */
  assign n1688_o = sndopc[4:0];
  /* TG68KdotC_Kernel.vhd:1307:67  */
  assign n1690_o = n1688_o - 5'b00001;
  /* TG68KdotC_Kernel.vhd:1304:17  */
  assign n1691_o = n1684_o ? n1687_o : n1690_o;
  /* TG68KdotC_Kernel.vhd:1309:37  */
  assign n1692_o = bf_width + bf_offset;
  /* TG68KdotC_Kernel.vhd:1310:43  */
  assign n1693_o = bf_bhits[3];
  /* TG68KdotC_Kernel.vhd:1310:31  */
  assign n1694_o = ~n1693_o;
  /* TG68KdotC_Kernel.vhd:1314:26  */
  assign n1695_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:1314:39  */
  assign n1697_o = n1695_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:1315:41  */
  assign n1699_o = 6'b100000 - bf_shift;
  assign n1702_o = n1699_o[4:0];
  assign n1703_o = bf_shift[4:0];
  /* TG68KdotC_Kernel.vhd:1314:17  */
  assign n1704_o = n1697_o ? n1702_o : n1703_o;
  /* TG68KdotC_Kernel.vhd:1321:26  */
  assign n1705_o = opcode[4:3];
  /* TG68KdotC_Kernel.vhd:1321:38  */
  assign n1707_o = n1705_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1322:34  */
  assign n1708_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:1322:47  */
  assign n1710_o = n1708_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:1323:53  */
  assign n1712_o = bf_bhits + 6'b000001;
  /* TG68KdotC_Kernel.vhd:1325:47  */
  assign n1714_o = 6'b011111 - bf_bhits;
  assign n1717_o = n1712_o[4:0];
  assign n1718_o = n1714_o[4:0];
  /* TG68KdotC_Kernel.vhd:1322:25  */
  assign n1719_o = n1710_o ? n1717_o : n1718_o;
  /* TG68KdotC_Kernel.vhd:1329:34  */
  assign n1720_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:1329:47  */
  assign n1722_o = n1720_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:1330:69  */
  assign n1723_o = bf_bhits[2:0];
  /* TG68KdotC_Kernel.vhd:1330:60  */
  assign n1725_o = {3'b000, n1723_o};
  /* TG68KdotC_Kernel.vhd:1330:53  */
  assign n1727_o = 6'b011001 + n1725_o;
  assign n1729_o = n1727_o[4:0];
  /* TG68KdotC_Kernel.vhd:1333:66  */
  assign n1730_o = bf_bhits[2:0];
  /* TG68KdotC_Kernel.vhd:1333:57  */
  assign n1732_o = 3'b111 - n1730_o;
  /* TG68KdotC_Kernel.vhd:1333:50  */
  assign n1734_o = {3'b000, n1732_o};
  assign n1735_o = {1'b0, n1729_o};
  /* TG68KdotC_Kernel.vhd:1329:25  */
  assign n1736_o = n1722_o ? n1735_o : n1734_o;
  assign n1738_o = n1672_o[4:3];
  assign n1739_o = n1675_o[4:3];
  /* TG68KdotC_Kernel.vhd:1291:17  */
  assign n1740_o = n1669_o ? n1738_o : n1739_o;
  /* TG68KdotC_Kernel.vhd:1321:17  */
  assign n1741_o = n1707_o ? n1740_o : 2'b00;
  assign n1742_o = n1672_o[5];
  assign n1743_o = n1675_o[5];
  /* TG68KdotC_Kernel.vhd:1291:17  */
  assign n1744_o = n1669_o ? n1742_o : n1743_o;
  assign n1745_o = n1672_o[2:0];
  assign n1746_o = n1675_o[2:0];
  /* TG68KdotC_Kernel.vhd:1291:17  */
  assign n1747_o = n1669_o ? n1745_o : n1746_o;
  assign n1748_o = {1'b0, n1719_o};
  /* TG68KdotC_Kernel.vhd:1321:17  */
  assign n1749_o = n1707_o ? n1748_o : n1736_o;
  /* TG68KdotC_Kernel.vhd:1338:30  */
  assign n1750_o = bf_bhits[5:3];
  /* TG68KdotC_Kernel.vhd:1339:25  */
  assign n1752_o = n1750_o == 3'b000;
  /* TG68KdotC_Kernel.vhd:1341:25  */
  assign n1754_o = n1750_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:1343:25  */
  assign n1756_o = n1750_o == 3'b010;
  /* TG68KdotC_Kernel.vhd:1345:25  */
  assign n1758_o = n1750_o == 3'b011;
  assign n1759_o = {n1758_o, n1756_o, n1754_o, n1752_o};
  /* TG68KdotC_Kernel.vhd:1338:17  */
  always @*
    case (n1759_o)
      4'b1000: n1765_o = 6'b100001;
      4'b0100: n1765_o = 6'b100011;
      4'b0010: n1765_o = 6'b100111;
      4'b0001: n1765_o = 6'b101111;
      default: n1765_o = 6'b100000;
    endcase
  /* TG68KdotC_Kernel.vhd:1350:28  */
  assign n1767_o = setstate == 2'b00;
  /* TG68KdotC_Kernel.vhd:1350:17  */
  assign n1769_o = n1767_o ? 6'b100111 : n1765_o;
  /* TG68KdotC_Kernel.vhd:1360:24  */
  assign n1773_o = exec[17];
  /* TG68KdotC_Kernel.vhd:1361:59  */
  assign n1774_o = last_data_read[15:8];
  /* TG68KdotC_Kernel.vhd:1361:41  */
  assign n1775_o = flagssr & n1774_o;
  /* TG68KdotC_Kernel.vhd:1362:27  */
  assign n1776_o = exec[18];
  /* TG68KdotC_Kernel.vhd:1363:59  */
  assign n1777_o = last_data_read[15:8];
  /* TG68KdotC_Kernel.vhd:1363:41  */
  assign n1778_o = flagssr ^ n1777_o;
  /* TG68KdotC_Kernel.vhd:1364:27  */
  assign n1779_o = exec[19];
  /* TG68KdotC_Kernel.vhd:1365:58  */
  assign n1780_o = last_data_read[15:8];
  /* TG68KdotC_Kernel.vhd:1365:41  */
  assign n1781_o = flagssr | n1780_o;
  /* TG68KdotC_Kernel.vhd:1367:39  */
  assign n1782_o = op2out[15:8];
  /* TG68KdotC_Kernel.vhd:1364:17  */
  assign n1783_o = n1779_o ? n1781_o : n1782_o;
  /* TG68KdotC_Kernel.vhd:1362:17  */
  assign n1784_o = n1776_o ? n1778_o : n1783_o;
  /* TG68KdotC_Kernel.vhd:1360:17  */
  assign n1785_o = n1773_o ? n1775_o : n1784_o;
  /* TG68KdotC_Kernel.vhd:1379:62  */
  assign n1788_o = flagssr[7];
  /* TG68KdotC_Kernel.vhd:1380:47  */
  assign n1789_o = set[41];
  /* TG68KdotC_Kernel.vhd:1381:59  */
  assign n1790_o = ~svmode;
  /* TG68KdotC_Kernel.vhd:1380:41  */
  assign n1791_o = n1789_o ? n1790_o : presvmode;
  /* TG68KdotC_Kernel.vhd:1378:33  */
  assign n1792_o = setopcode ? n1788_o : make_trace;
  /* TG68KdotC_Kernel.vhd:1377:25  */
  assign n1793_o = n1880_o ? n1791_o : svmode;
  /* TG68KdotC_Kernel.vhd:1386:50  */
  assign n1794_o = trap_berr | trap_illegal;
  /* TG68KdotC_Kernel.vhd:1386:70  */
  assign n1795_o = n1794_o | trap_addr_error;
  /* TG68KdotC_Kernel.vhd:1386:93  */
  assign n1796_o = n1795_o | trap_priv;
  /* TG68KdotC_Kernel.vhd:1386:110  */
  assign n1797_o = n1796_o | trap_1010;
  /* TG68KdotC_Kernel.vhd:1386:127  */
  assign n1798_o = n1797_o | trap_1111;
  assign n1800_o = flagssr[7];
  /* TG68KdotC_Kernel.vhd:1386:33  */
  assign n1801_o = n1798_o ? 1'b0 : n1800_o;
  /* TG68KdotC_Kernel.vhd:1386:33  */
  assign n1803_o = n1798_o ? 1'b0 : n1792_o;
  /* TG68KdotC_Kernel.vhd:1390:39  */
  assign n1804_o = set[41];
  /* TG68KdotC_Kernel.vhd:1391:54  */
  assign n1805_o = ~presvmode;
  /* TG68KdotC_Kernel.vhd:1392:55  */
  assign n1806_o = ~presvmode;
  /* TG68KdotC_Kernel.vhd:1393:50  */
  assign n1807_o = ~presvmode;
  assign n1808_o = n9781_o[2];
  /* TG68KdotC_Kernel.vhd:1390:33  */
  assign n1809_o = n1804_o ? n1807_o : n1808_o;
  assign n1810_o = flagssr[5];
  /* TG68KdotC_Kernel.vhd:1390:33  */
  assign n1811_o = n1804_o ? n1806_o : n1810_o;
  /* TG68KdotC_Kernel.vhd:1377:25  */
  assign n1812_o = n1881_o ? n1805_o : presvmode;
  /* TG68KdotC_Kernel.vhd:1395:47  */
  assign n1814_o = micro_state == 7'b0110110;
  /* TG68KdotC_Kernel.vhd:1395:33  */
  assign n1816_o = n1814_o ? 1'b0 : n1801_o;
  /* TG68KdotC_Kernel.vhd:1398:60  */
  assign n1818_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:1398:51  */
  assign n1819_o = n1818_o & trap_trace;
  /* TG68KdotC_Kernel.vhd:1398:33  */
  assign n1821_o = n1819_o ? 1'b0 : n1803_o;
  /* TG68KdotC_Kernel.vhd:1401:40  */
  assign n1822_o = exec[59];
  /* TG68KdotC_Kernel.vhd:1401:55  */
  assign n1823_o = n1822_o | set_stop;
  assign n1825_o = flagssr[4:0];
  assign n1826_o = flagssr[6];
  assign n1827_o = {n1816_o, n1826_o, n1811_o, n1825_o};
  /* TG68KdotC_Kernel.vhd:1404:50  */
  assign n1829_o = trap_interrupt & interrupt;
  assign n1830_o = data_read[10:8];
  assign n1831_o = n1827_o[2:0];
  /* TG68KdotC_Kernel.vhd:1401:33  */
  assign n1832_o = n1823_o ? n1830_o : n1831_o;
  /* TG68KdotC_Kernel.vhd:1404:33  */
  assign n1833_o = n1829_o ? ripl_nr : n1832_o;
  assign n1834_o = data_read[15:11];
  assign n1835_o = n1827_o[7:3];
  /* TG68KdotC_Kernel.vhd:1401:33  */
  assign n1836_o = n1823_o ? n1834_o : n1835_o;
  /* TG68KdotC_Kernel.vhd:1407:40  */
  assign n1837_o = exec[52];
  /* TG68KdotC_Kernel.vhd:1409:54  */
  assign n1838_o = srin[5];
  /* TG68KdotC_Kernel.vhd:1410:43  */
  assign n1839_o = exec[35];
  /* TG68KdotC_Kernel.vhd:1411:57  */
  assign n1840_o = flagssr[5];
  /* TG68KdotC_Kernel.vhd:1410:33  */
  assign n1841_o = n1839_o ? n1840_o : n1809_o;
  /* TG68KdotC_Kernel.vhd:1407:33  */
  assign n1842_o = n1837_o ? n1838_o : n1841_o;
  assign n1843_o = {n1836_o, n1833_o};
  /* TG68KdotC_Kernel.vhd:1413:33  */
  assign n1846_o = interrupt ? 1'b1 : n1842_o;
  /* TG68KdotC_Kernel.vhd:1416:39  */
  assign n1847_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:1416:42  */
  assign n1848_o = ~n1847_o;
  assign n1851_o = srin[4];
  assign n1852_o = n1843_o[4];
  /* TG68KdotC_Kernel.vhd:1407:33  */
  assign n1853_o = n1837_o ? n1851_o : n1852_o;
  /* TG68KdotC_Kernel.vhd:1416:33  */
  assign n1854_o = n1848_o ? 1'b0 : n1853_o;
  assign n1855_o = srin[6];
  assign n1856_o = n1843_o[6];
  /* TG68KdotC_Kernel.vhd:1407:33  */
  assign n1857_o = n1837_o ? n1855_o : n1856_o;
  /* TG68KdotC_Kernel.vhd:1416:33  */
  assign n1858_o = n1848_o ? 1'b0 : n1857_o;
  assign n1865_o = srin[7];
  assign n1866_o = n1843_o[7];
  /* TG68KdotC_Kernel.vhd:1407:33  */
  assign n1867_o = n1837_o ? n1865_o : n1866_o;
  assign n1868_o = srin[5];
  assign n1869_o = n1843_o[5];
  /* TG68KdotC_Kernel.vhd:1407:33  */
  assign n1870_o = n1837_o ? n1868_o : n1869_o;
  assign n1872_o = srin[2:0];
  assign n1873_o = n1843_o[2:0];
  /* TG68KdotC_Kernel.vhd:1407:33  */
  assign n1874_o = n1837_o ? n1872_o : n1873_o;
  assign n1875_o = n9781_o[2];
  /* TG68KdotC_Kernel.vhd:1377:25  */
  assign n1876_o = clkena_lw ? n1846_o : n1875_o;
  assign n1877_o = {n1867_o, n1858_o, n1870_o, n1854_o, 1'b0, n1874_o};
  /* TG68KdotC_Kernel.vhd:1377:25  */
  assign n1878_o = clkena_lw ? n1877_o : flagssr;
  /* TG68KdotC_Kernel.vhd:1377:25  */
  assign n1879_o = clkena_lw ? n1821_o : make_trace;
  /* TG68KdotC_Kernel.vhd:1377:25  */
  assign n1880_o = setopcode & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1377:25  */
  assign n1881_o = n1804_o & clkena_lw;
  /* TG68KdotC_Kernel.vhd:1371:25  */
  assign n1882_o = reset ? 1'b1 : n1876_o;
  /* TG68KdotC_Kernel.vhd:1371:25  */
  assign n1884_o = reset ? 8'b00100111 : n1878_o;
  /* TG68KdotC_Kernel.vhd:1371:25  */
  assign n1886_o = reset ? 1'b0 : n1879_o;
  /* TG68KdotC_Kernel.vhd:1371:25  */
  assign n1888_o = reset ? 1'b1 : n1793_o;
  /* TG68KdotC_Kernel.vhd:1371:25  */
  assign n1890_o = reset ? 1'b1 : n1812_o;
  /* TG68KdotC_Kernel.vhd:1453:39  */
  assign n1900_o = opcode[4:3];
  /* TG68KdotC_Kernel.vhd:1495:27  */
  assign n1902_o = rot_cnt != 6'b000001;
  /* TG68KdotC_Kernel.vhd:1496:47  */
  assign n1904_o = rot_cnt - 6'b000001;
  /* TG68KdotC_Kernel.vhd:1495:17  */
  assign n1906_o = n1902_o ? n1904_o : 6'b000001;
  /* TG68KdotC_Kernel.vhd:1507:28  */
  assign n1912_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:1508:25  */
  assign n1914_o = n1912_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1509:25  */
  assign n1916_o = n1912_o == 2'b01;
  assign n1917_o = {n1916_o, n1914_o};
  /* TG68KdotC_Kernel.vhd:1507:17  */
  always @*
    case (n1917_o)
      2'b10: n1921_o = 2'b01;
      2'b01: n1921_o = 2'b00;
      default: n1921_o = 2'b10;
    endcase
  /* TG68KdotC_Kernel.vhd:1513:32  */
  assign n1922_o = exec_write_back & execopc;
  assign n1924_o = n1909_o[83];
  /* TG68KdotC_Kernel.vhd:1513:17  */
  assign n1925_o = n1922_o ? 1'b1 : n1924_o;
  /* TG68KdotC_Kernel.vhd:1517:34  */
  assign n1928_o = trap_berr & interrupt;
  /* TG68KdotC_Kernel.vhd:1519:37  */
  assign n1929_o = ~presvmode;
  assign n1931_o = n1909_o[41];
  /* TG68KdotC_Kernel.vhd:1517:17  */
  assign n1932_o = n1938_o ? 1'b1 : n1931_o;
  /* TG68KdotC_Kernel.vhd:1517:17  */
  assign n1935_o = n1928_o ? 2'b01 : 2'b00;
  /* TG68KdotC_Kernel.vhd:1517:17  */
  assign n1938_o = n1929_o & n1928_o;
  assign n1940_o = n1909_o[40:39];
  /* TG68KdotC_Kernel.vhd:1517:17  */
  assign n1943_o = n1928_o ? 7'b0110111 : 7'b0000000;
  /* TG68KdotC_Kernel.vhd:1524:42  */
  assign n1945_o = ~trapd;
  /* TG68KdotC_Kernel.vhd:1524:33  */
  assign n1946_o = n1945_o & trapmake;
  /* TG68KdotC_Kernel.vhd:1525:31  */
  assign n1947_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:1525:59  */
  assign n1948_o = trap_trapv | set_z_error;
  /* TG68KdotC_Kernel.vhd:1525:85  */
  assign n1949_o = exec[43];
  /* TG68KdotC_Kernel.vhd:1525:78  */
  assign n1950_o = n1948_o | n1949_o;
  /* TG68KdotC_Kernel.vhd:1525:39  */
  assign n1951_o = n1950_o & n1947_o;
  /* TG68KdotC_Kernel.vhd:1527:25  */
  assign n1954_o = trap_addr_error ? 7'b0110111 : 7'b0110011;
  /* TG68KdotC_Kernel.vhd:1525:25  */
  assign n1956_o = n1951_o ? 7'b0110010 : n1954_o;
  /* TG68KdotC_Kernel.vhd:1532:46  */
  assign n1957_o = ~use_vbr_stackframe;
  assign n1959_o = n1909_o[25];
  /* TG68KdotC_Kernel.vhd:1524:17  */
  assign n1960_o = n1967_o ? 1'b1 : n1959_o;
  /* TG68KdotC_Kernel.vhd:1536:37  */
  assign n1961_o = ~presvmode;
  /* TG68KdotC_Kernel.vhd:1524:17  */
  assign n1963_o = n1968_o ? 1'b1 : n1932_o;
  /* TG68KdotC_Kernel.vhd:1524:17  */
  assign n1965_o = n1946_o ? 2'b01 : n1935_o;
  /* TG68KdotC_Kernel.vhd:1524:17  */
  assign n1967_o = n1957_o & n1946_o;
  /* TG68KdotC_Kernel.vhd:1524:17  */
  assign n1968_o = n1961_o & n1946_o;
  /* TG68KdotC_Kernel.vhd:1524:17  */
  assign n1971_o = n1946_o ? n1956_o : n1943_o;
  /* TG68KdotC_Kernel.vhd:1541:31  */
  assign n1973_o = micro_state == 7'b0100111;
  /* TG68KdotC_Kernel.vhd:1541:55  */
  assign n1974_o = trap_trace & interrupt;
  /* TG68KdotC_Kernel.vhd:1541:37  */
  assign n1975_o = n1973_o | n1974_o;
  /* TG68KdotC_Kernel.vhd:1543:50  */
  assign n1976_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:1543:43  */
  assign n1977_o = n1976_o & trap_trace;
  /* TG68KdotC_Kernel.vhd:1543:25  */
  assign n1980_o = n1977_o ? 7'b0110010 : 7'b0110011;
  /* TG68KdotC_Kernel.vhd:1553:37  */
  assign n1981_o = ~presvmode;
  /* TG68KdotC_Kernel.vhd:1541:17  */
  assign n1983_o = n1986_o ? 1'b1 : n1963_o;
  /* TG68KdotC_Kernel.vhd:1541:17  */
  assign n1985_o = n1975_o ? 2'b01 : n1965_o;
  /* TG68KdotC_Kernel.vhd:1541:17  */
  assign n1986_o = n1981_o & n1975_o;
  /* TG68KdotC_Kernel.vhd:1541:17  */
  assign n1987_o = n1975_o ? n1980_o : n1971_o;
  /* TG68KdotC_Kernel.vhd:1558:24  */
  assign n1989_o = micro_state == 7'b0100111;
  /* TG68KdotC_Kernel.vhd:1558:51  */
  assign n1990_o = trap_trace & interrupt;
  /* TG68KdotC_Kernel.vhd:1558:31  */
  assign n1991_o = n1989_o | n1990_o;
  /* TG68KdotC_Kernel.vhd:1559:24  */
  assign n1992_o = ~presvmode;
  /* TG68KdotC_Kernel.vhd:1558:9  */
  assign n1994_o = n1997_o ? 1'b1 : n1983_o;
  /* TG68KdotC_Kernel.vhd:1558:9  */
  assign n1996_o = n1991_o ? 2'b01 : n1985_o;
  /* TG68KdotC_Kernel.vhd:1558:9  */
  assign n1997_o = n1992_o & n1991_o;
  /* TG68KdotC_Kernel.vhd:1565:46  */
  assign n1998_o = flagssr[5];
  /* TG68KdotC_Kernel.vhd:1565:49  */
  assign n1999_o = n1998_o != presvmode;
  /* TG68KdotC_Kernel.vhd:1565:35  */
  assign n2000_o = n1999_o & setexecopc;
  /* TG68KdotC_Kernel.vhd:1565:17  */
  assign n2002_o = n2000_o ? 1'b1 : n1994_o;
  /* TG68KdotC_Kernel.vhd:1571:34  */
  assign n2003_o = trap_interrupt & interrupt;
  /* TG68KdotC_Kernel.vhd:1571:17  */
  assign n2006_o = n2003_o ? 2'b10 : n1996_o;
  /* TG68KdotC_Kernel.vhd:1571:17  */
  assign n2007_o = n2003_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1571:17  */
  assign n2009_o = n2003_o ? 7'b0100111 : n1987_o;
  /* TG68KdotC_Kernel.vhd:1578:23  */
  assign n2010_o = set[41];
  /* TG68KdotC_Kernel.vhd:1578:17  */
  assign n2015_o = n2010_o ? 1'b1 : 1'b0;
  assign n2017_o = {1'b1, 1'b1};
  assign n2018_o = n1909_o[66:65];
  /* TG68KdotC_Kernel.vhd:1578:17  */
  assign n2019_o = n2010_o ? n2017_o : n2018_o;
  /* TG68KdotC_Kernel.vhd:1584:27  */
  assign n2022_o = ~ea_only;
  /* TG68KdotC_Kernel.vhd:1584:39  */
  assign n2023_o = set[62];
  /* TG68KdotC_Kernel.vhd:1584:32  */
  assign n2024_o = n2023_o & n2022_o;
  /* TG68KdotC_Kernel.vhd:1584:17  */
  assign n2026_o = n2024_o ? 2'b10 : n2006_o;
  /* TG68KdotC_Kernel.vhd:1590:28  */
  assign n2027_o = setstate[1];
  /* TG68KdotC_Kernel.vhd:1590:52  */
  assign n2028_o = set_datatype[1];
  /* TG68KdotC_Kernel.vhd:1590:36  */
  assign n2029_o = n2028_o & n2027_o;
  assign n2031_o = n1909_o[73];
  /* TG68KdotC_Kernel.vhd:1590:17  */
  assign n2032_o = n2029_o ? 1'b1 : n2031_o;
  /* TG68KdotC_Kernel.vhd:1594:38  */
  assign n2035_o = decodeopc & ea_build_now;
  /* TG68KdotC_Kernel.vhd:1594:64  */
  assign n2036_o = exec[42];
  /* TG68KdotC_Kernel.vhd:1594:57  */
  assign n2037_o = n2035_o | n2036_o;
  /* TG68KdotC_Kernel.vhd:1595:36  */
  assign n2038_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1599:50  */
  assign n2040_o = opcode[3];
  /* TG68KdotC_Kernel.vhd:1601:58  */
  assign n2042_o = opcode[2:0];
  /* TG68KdotC_Kernel.vhd:1601:70  */
  assign n2044_o = n2042_o == 3'b111;
  assign n2046_o = n1909_o[50];
  /* TG68KdotC_Kernel.vhd:1599:41  */
  assign n2047_o = n2051_o ? 1'b1 : n2046_o;
  assign n2048_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1599:41  */
  assign n2049_o = n2040_o ? 1'b1 : n2048_o;
  /* TG68KdotC_Kernel.vhd:1599:41  */
  assign n2051_o = n2044_o & n2040_o;
  /* TG68KdotC_Kernel.vhd:1605:50  */
  assign n2052_o = opcode[5];
  /* TG68KdotC_Kernel.vhd:1607:58  */
  assign n2054_o = opcode[2:0];
  /* TG68KdotC_Kernel.vhd:1607:70  */
  assign n2056_o = n2054_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:1605:41  */
  assign n2058_o = n2061_o ? 1'b1 : n2047_o;
  assign n2059_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1605:41  */
  assign n2060_o = n2052_o ? 1'b1 : n2059_o;
  /* TG68KdotC_Kernel.vhd:1605:41  */
  assign n2061_o = n2056_o & n2052_o;
  /* TG68KdotC_Kernel.vhd:1596:33  */
  assign n2063_o = n2038_o == 3'b010;
  /* TG68KdotC_Kernel.vhd:1596:43  */
  assign n2065_o = n2038_o == 3'b011;
  /* TG68KdotC_Kernel.vhd:1596:43  */
  assign n2066_o = n2063_o | n2065_o;
  /* TG68KdotC_Kernel.vhd:1596:49  */
  assign n2068_o = n2038_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:1596:49  */
  assign n2069_o = n2066_o | n2068_o;
  /* TG68KdotC_Kernel.vhd:1611:33  */
  assign n2071_o = n2038_o == 3'b101;
  /* TG68KdotC_Kernel.vhd:1613:33  */
  assign n2073_o = n2038_o == 3'b110;
  /* TG68KdotC_Kernel.vhd:1617:52  */
  assign n2074_o = opcode[2:0];
  /* TG68KdotC_Kernel.vhd:1618:49  */
  assign n2076_o = n2074_o == 3'b000;
  /* TG68KdotC_Kernel.vhd:1620:49  */
  assign n2079_o = n2074_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:1623:49  */
  assign n2082_o = n2074_o == 3'b010;
  /* TG68KdotC_Kernel.vhd:1628:49  */
  assign n2085_o = n2074_o == 3'b011;
  /* TG68KdotC_Kernel.vhd:1637:68  */
  assign n2087_o = datatype == 2'b10;
  /* TG68KdotC_Kernel.vhd:1637:57  */
  assign n2089_o = n2087_o ? 1'b1 : n2032_o;
  /* TG68KdotC_Kernel.vhd:1634:49  */
  assign n2091_o = n2074_o == 3'b100;
  assign n2092_o = {n2091_o, n2085_o, n2082_o, n2079_o, n2076_o};
  /* TG68KdotC_Kernel.vhd:1617:41  */
  always @*
    case (n2092_o)
      5'b10000: n2095_o = 1'b1;
      5'b01000: n2095_o = 1'b0;
      5'b00100: n2095_o = 1'b0;
      5'b00010: n2095_o = 1'b0;
      5'b00001: n2095_o = 1'b0;
      default: n2095_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1617:41  */
  always @*
    case (n2092_o)
      5'b10000: n2098_o = 1'b0;
      5'b01000: n2098_o = 1'b1;
      5'b00100: n2098_o = 1'b0;
      5'b00010: n2098_o = 1'b0;
      5'b00001: n2098_o = 1'b0;
      default: n2098_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1617:41  */
  always @*
    case (n2092_o)
      5'b10000: n2101_o = 1'b1;
      5'b01000: n2101_o = 1'b0;
      5'b00100: n2101_o = 1'b0;
      5'b00010: n2101_o = 1'b0;
      5'b00001: n2101_o = 1'b0;
      default: n2101_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1617:41  */
  always @*
    case (n2092_o)
      5'b10000: n2105_o = 1'b0;
      5'b01000: n2105_o = 1'b1;
      5'b00100: n2105_o = 1'b1;
      5'b00010: n2105_o = 1'b0;
      5'b00001: n2105_o = 1'b0;
      default: n2105_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1617:41  */
  always @*
    case (n2092_o)
      5'b10000: n2109_o = 1'b0;
      5'b01000: n2109_o = 1'b1;
      5'b00100: n2109_o = 1'b1;
      5'b00010: n2109_o = 1'b0;
      5'b00001: n2109_o = 1'b0;
      default: n2109_o = 1'b0;
    endcase
  assign n2110_o = n1909_o[22];
  /* TG68KdotC_Kernel.vhd:1617:41  */
  always @*
    case (n2092_o)
      5'b10000: n2111_o = n2110_o;
      5'b01000: n2111_o = 1'b1;
      5'b00100: n2111_o = 1'b1;
      5'b00010: n2111_o = n2110_o;
      5'b00001: n2111_o = n2110_o;
      default: n2111_o = n2110_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1617:41  */
  always @*
    case (n2092_o)
      5'b10000: n2112_o = n2089_o;
      5'b01000: n2112_o = n2032_o;
      5'b00100: n2112_o = n2032_o;
      5'b00010: n2112_o = 1'b1;
      5'b00001: n2112_o = n2032_o;
      default: n2112_o = n2032_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1617:41  */
  always @*
    case (n2092_o)
      5'b10000: n2117_o = n2009_o;
      5'b01000: n2117_o = 7'b0000101;
      5'b00100: n2117_o = 7'b0000100;
      5'b00010: n2117_o = 7'b0000010;
      5'b00001: n2117_o = 7'b0000010;
      default: n2117_o = n2009_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1616:33  */
  assign n2119_o = n2038_o == 3'b111;
  assign n2120_o = {n2119_o, n2073_o, n2071_o, n2069_o};
  /* TG68KdotC_Kernel.vhd:1595:25  */
  always @*
    case (n2120_o)
      4'b1000: n2123_o = n2095_o;
      4'b0100: n2123_o = 1'b0;
      4'b0010: n2123_o = 1'b0;
      4'b0001: n2123_o = 1'b1;
      default: n2123_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1595:25  */
  always @*
    case (n2120_o)
      4'b1000: n2126_o = n2098_o;
      4'b0100: n2126_o = 1'b1;
      4'b0010: n2126_o = 1'b0;
      4'b0001: n2126_o = 1'b0;
      default: n2126_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1595:25  */
  always @*
    case (n2120_o)
      4'b1000: n2128_o = n2101_o;
      4'b0100: n2128_o = 1'b0;
      4'b0010: n2128_o = 1'b0;
      4'b0001: n2128_o = 1'b0;
      default: n2128_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1595:25  */
  always @*
    case (n2120_o)
      4'b1000: n2130_o = n2105_o;
      4'b0100: n2130_o = 1'b0;
      4'b0010: n2130_o = 1'b0;
      4'b0001: n2130_o = 1'b0;
      default: n2130_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1595:25  */
  always @*
    case (n2120_o)
      4'b1000: n2132_o = n2109_o;
      4'b0100: n2132_o = 1'b0;
      4'b0010: n2132_o = 1'b0;
      4'b0001: n2132_o = 1'b0;
      default: n2132_o = 1'b0;
    endcase
  assign n2133_o = n1909_o[22];
  /* TG68KdotC_Kernel.vhd:1595:25  */
  always @*
    case (n2120_o)
      4'b1000: n2134_o = n2111_o;
      4'b0100: n2134_o = n2133_o;
      4'b0010: n2134_o = n2133_o;
      4'b0001: n2134_o = n2133_o;
      default: n2134_o = n2133_o;
    endcase
  assign n2135_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1595:25  */
  always @*
    case (n2120_o)
      4'b1000: n2136_o = n2135_o;
      4'b0100: n2136_o = n2135_o;
      4'b0010: n2136_o = n2135_o;
      4'b0001: n2136_o = n2049_o;
      default: n2136_o = n2135_o;
    endcase
  assign n2137_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1595:25  */
  always @*
    case (n2120_o)
      4'b1000: n2138_o = n2137_o;
      4'b0100: n2138_o = n2137_o;
      4'b0010: n2138_o = n2137_o;
      4'b0001: n2138_o = n2060_o;
      default: n2138_o = n2137_o;
    endcase
  assign n2139_o = n1909_o[50];
  /* TG68KdotC_Kernel.vhd:1595:25  */
  always @*
    case (n2120_o)
      4'b1000: n2140_o = n2139_o;
      4'b0100: n2140_o = n2139_o;
      4'b0010: n2140_o = n2139_o;
      4'b0001: n2140_o = n2058_o;
      default: n2140_o = n2139_o;
    endcase
  assign n2141_o = n1909_o[62];
  /* TG68KdotC_Kernel.vhd:1595:25  */
  always @*
    case (n2120_o)
      4'b1000: n2142_o = n2141_o;
      4'b0100: n2142_o = n2141_o;
      4'b0010: n2142_o = n2141_o;
      4'b0001: n2142_o = 1'b1;
      default: n2142_o = n2141_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1595:25  */
  always @*
    case (n2120_o)
      4'b1000: n2143_o = n2112_o;
      4'b0100: n2143_o = n2032_o;
      4'b0010: n2143_o = n2032_o;
      4'b0001: n2143_o = n2032_o;
      default: n2143_o = n2032_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1595:25  */
  always @*
    case (n2120_o)
      4'b1000: n2146_o = n2117_o;
      4'b0100: n2146_o = 7'b0000101;
      4'b0010: n2146_o = 7'b0000100;
      4'b0001: n2146_o = n2009_o;
      default: n2146_o = n2009_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n2148_o = n2037_o ? n2123_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n2151_o = n2037_o ? n2126_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n2154_o = n2037_o ? n2128_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n2157_o = n2037_o ? n2130_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n2160_o = n2037_o ? n2132_o : 1'b0;
  assign n2162_o = {n2138_o, n2136_o};
  assign n2163_o = n1909_o[22];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n2164_o = n2037_o ? n2134_o : n2163_o;
  assign n2165_o = n1909_o[47:46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n2166_o = n2037_o ? n2162_o : n2165_o;
  assign n2167_o = n1909_o[50];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n2168_o = n2037_o ? n2140_o : n2167_o;
  assign n2169_o = n1909_o[62];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n2170_o = n2037_o ? n2142_o : n2169_o;
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n2171_o = n2037_o ? n2143_o : n2032_o;
  assign n2177_o = n1909_o[49:48];
  assign n2178_o = n1909_o[64:63];
  assign n2179_o = n1909_o[61:51];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n2180_o = n2037_o ? n2146_o : n2009_o;
  /* TG68KdotC_Kernel.vhd:1649:28  */
  assign n2181_o = tg68_pc[0];
  /* TG68KdotC_Kernel.vhd:1649:54  */
  assign n2183_o = micro_state == 7'b0000001;
  /* TG68KdotC_Kernel.vhd:1649:38  */
  assign n2184_o = n2183_o & n2181_o;
  /* TG68KdotC_Kernel.vhd:1653:28  */
  assign n2185_o = opcode[15:12];
  /* TG68KdotC_Kernel.vhd:1656:34  */
  assign n2186_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:1656:52  */
  assign n2187_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1656:64  */
  assign n2189_o = n2187_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:1656:42  */
  assign n2190_o = n2189_o & n2186_o;
  /* TG68KdotC_Kernel.vhd:1660:42  */
  assign n2193_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:1660:45  */
  assign n2194_o = ~n2193_o;
  assign n2198_o = n1909_o[37];
  /* TG68KdotC_Kernel.vhd:1660:33  */
  assign n2199_o = n2194_o ? 1'b1 : n2198_o;
  /* TG68KdotC_Kernel.vhd:1660:33  */
  assign n2201_o = n2194_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1660:33  */
  assign n2203_o = n2194_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1666:50  */
  assign n2204_o = opcode[6];
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2206_o = n2212_o ? 1'b1 : n2199_o;
  /* TG68KdotC_Kernel.vhd:1669:50  */
  assign n2207_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:1669:53  */
  assign n2208_o = ~n2207_o;
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2210_o = n2211_o ? 1'b1 : n2154_o;
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2211_o = n2208_o & decodeopc;
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2212_o = n2204_o & decodeopc;
  /* TG68KdotC_Kernel.vhd:1665:33  */
  assign n2214_o = decodeopc ? 7'b1001110 : n2180_o;
  /* TG68KdotC_Kernel.vhd:1674:33  */
  assign n2217_o = setexecopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1678:42  */
  assign n2218_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:1678:59  */
  assign n2219_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:1678:72  */
  assign n2221_o = n2219_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:1678:50  */
  assign n2222_o = n2218_o | n2221_o;
  /* TG68KdotC_Kernel.vhd:1679:50  */
  assign n2223_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1679:62  */
  assign n2225_o = n2223_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:1680:51  */
  assign n2226_o = opcode[8:3];
  /* TG68KdotC_Kernel.vhd:1680:63  */
  assign n2228_o = n2226_o != 6'b000111;
  /* TG68KdotC_Kernel.vhd:1680:83  */
  assign n2229_o = opcode[2];
  /* TG68KdotC_Kernel.vhd:1680:86  */
  assign n2230_o = ~n2229_o;
  /* TG68KdotC_Kernel.vhd:1680:74  */
  assign n2231_o = n2228_o | n2230_o;
  /* TG68KdotC_Kernel.vhd:1679:70  */
  assign n2232_o = n2231_o & n2225_o;
  /* TG68KdotC_Kernel.vhd:1681:51  */
  assign n2233_o = opcode[8:2];
  /* TG68KdotC_Kernel.vhd:1681:63  */
  assign n2235_o = n2233_o != 7'b1001111;
  /* TG68KdotC_Kernel.vhd:1681:84  */
  assign n2236_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:1681:96  */
  assign n2238_o = n2236_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1681:75  */
  assign n2239_o = n2235_o | n2238_o;
  /* TG68KdotC_Kernel.vhd:1680:92  */
  assign n2240_o = n2239_o & n2232_o;
  /* TG68KdotC_Kernel.vhd:1682:51  */
  assign n2241_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:1682:63  */
  assign n2243_o = n2241_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1682:78  */
  assign n2244_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1682:90  */
  assign n2246_o = n2244_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:1682:69  */
  assign n2247_o = n2243_o | n2246_o;
  /* TG68KdotC_Kernel.vhd:1682:107  */
  assign n2248_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:1682:119  */
  assign n2250_o = n2248_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1682:98  */
  assign n2251_o = n2247_o | n2250_o;
  /* TG68KdotC_Kernel.vhd:1681:103  */
  assign n2252_o = n2251_o & n2240_o;
  /* TG68KdotC_Kernel.vhd:1685:58  */
  assign n2255_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:1685:70  */
  assign n2257_o = n2255_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:1686:66  */
  assign n2258_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:1686:78  */
  assign n2260_o = n2258_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1686:57  */
  assign n2263_o = n2260_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1685:49  */
  assign n2266_o = n2257_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1685:49  */
  assign n2268_o = n2257_o ? n2263_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1691:58  */
  assign n2269_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:1691:70  */
  assign n2271_o = n2269_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1691:49  */
  assign n2274_o = n2271_o ? 2'b10 : 2'b00;
  /* TG68KdotC_Kernel.vhd:1696:58  */
  assign n2275_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:1696:61  */
  assign n2276_o = ~n2275_o;
  assign n2279_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:1679:41  */
  assign n2280_o = n2305_o ? 1'b1 : n2279_o;
  assign n2281_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:1679:41  */
  assign n2282_o = n2307_o ? 1'b1 : n2281_o;
  /* TG68KdotC_Kernel.vhd:1679:41  */
  assign n2284_o = n2314_o ? 7'b0000001 : n2180_o;
  /* TG68KdotC_Kernel.vhd:1696:49  */
  assign n2287_o = n2276_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1696:49  */
  assign n2289_o = decodeopc & n2276_o;
  /* TG68KdotC_Kernel.vhd:1696:49  */
  assign n2291_o = decodeopc & n2276_o;
  /* TG68KdotC_Kernel.vhd:1696:49  */
  assign n2292_o = decodeopc & n2276_o;
  /* TG68KdotC_Kernel.vhd:1679:41  */
  assign n2293_o = n2252_o ? n2274_o : n1921_o;
  /* TG68KdotC_Kernel.vhd:1679:41  */
  assign n2295_o = n2252_o ? n2266_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1679:41  */
  assign n2298_o = n2252_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1679:41  */
  assign n2301_o = n2252_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1679:41  */
  assign n2303_o = n2252_o ? n2287_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1679:41  */
  assign n2305_o = n2289_o & n2252_o;
  /* TG68KdotC_Kernel.vhd:1679:41  */
  assign n2307_o = n2291_o & n2252_o;
  /* TG68KdotC_Kernel.vhd:1679:41  */
  assign n2309_o = n2252_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1679:41  */
  assign n2311_o = n2252_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1679:41  */
  assign n2313_o = n2252_o ? n2268_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1679:41  */
  assign n2314_o = n2292_o & n2252_o;
  /* TG68KdotC_Kernel.vhd:1709:45  */
  assign n2315_o = opcode[8:6];
  /* TG68KdotC_Kernel.vhd:1709:57  */
  assign n2317_o = n2315_o == 3'b011;
  /* TG68KdotC_Kernel.vhd:1710:47  */
  assign n2318_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:1711:58  */
  assign n2319_o = opcode[11];
  /* TG68KdotC_Kernel.vhd:1712:67  */
  assign n2320_o = opcode[10:9];
  /* TG68KdotC_Kernel.vhd:1712:80  */
  assign n2322_o = n2320_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:1713:66  */
  assign n2323_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:1713:78  */
  assign n2325_o = n2323_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:1712:87  */
  assign n2326_o = n2325_o & n2322_o;
  /* TG68KdotC_Kernel.vhd:1713:96  */
  assign n2327_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1713:108  */
  assign n2329_o = n2327_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:1713:125  */
  assign n2330_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:1713:137  */
  assign n2332_o = n2330_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1713:116  */
  assign n2333_o = n2329_o | n2332_o;
  /* TG68KdotC_Kernel.vhd:1713:85  */
  assign n2334_o = n2333_o & n2326_o;
  /* TG68KdotC_Kernel.vhd:1714:67  */
  assign n2335_o = opcode[10];
  /* TG68KdotC_Kernel.vhd:1714:86  */
  assign n2336_o = opcode[5:0];
  /* TG68KdotC_Kernel.vhd:1714:98  */
  assign n2338_o = n2336_o == 6'b111100;
  /* TG68KdotC_Kernel.vhd:1714:76  */
  assign n2339_o = n2338_o & n2335_o;
  /* TG68KdotC_Kernel.vhd:1713:145  */
  assign n2340_o = n2334_o | n2339_o;
  /* TG68KdotC_Kernel.vhd:1715:76  */
  assign n2341_o = opcode[10:9];
  /* TG68KdotC_Kernel.vhd:1716:73  */
  assign n2343_o = n2341_o == 2'b01;
  /* TG68KdotC_Kernel.vhd:1717:73  */
  assign n2345_o = n2341_o == 2'b10;
  assign n2346_o = {n2345_o, n2343_o};
  /* TG68KdotC_Kernel.vhd:1715:65  */
  always @*
    case (n2346_o)
      2'b10: n2350_o = 2'b01;
      2'b01: n2350_o = 2'b00;
      default: n2350_o = 2'b10;
    endcase
  /* TG68KdotC_Kernel.vhd:1720:74  */
  assign n2351_o = opcode[10];
  /* TG68KdotC_Kernel.vhd:1720:93  */
  assign n2352_o = opcode[5:0];
  /* TG68KdotC_Kernel.vhd:1720:105  */
  assign n2354_o = n2352_o == 6'b111100;
  /* TG68KdotC_Kernel.vhd:1720:83  */
  assign n2355_o = n2354_o & n2351_o;
  assign n2357_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:1721:73  */
  assign n2358_o = decodeopc ? 1'b1 : n2357_o;
  /* TG68KdotC_Kernel.vhd:1721:73  */
  assign n2360_o = decodeopc ? 7'b1000000 : n2180_o;
  assign n2363_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:1726:73  */
  assign n2364_o = decodeopc ? 1'b1 : n2363_o;
  assign n2365_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:1726:73  */
  assign n2366_o = decodeopc ? 1'b1 : n2365_o;
  /* TG68KdotC_Kernel.vhd:1726:73  */
  assign n2368_o = decodeopc ? 7'b0000001 : n2180_o;
  /* TG68KdotC_Kernel.vhd:1731:87  */
  assign n2370_o = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:1731:93  */
  assign n2371_o = nextpass & n2370_o;
  /* TG68KdotC_Kernel.vhd:1731:73  */
  assign n2377_o = n2371_o ? 2'b01 : n2026_o;
  /* TG68KdotC_Kernel.vhd:1731:73  */
  assign n2380_o = n2371_o ? 1'b1 : 1'b0;
  assign n2381_o = n1909_o[26];
  /* TG68KdotC_Kernel.vhd:1731:73  */
  assign n2382_o = n2371_o ? 1'b1 : n2381_o;
  assign n2383_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:1731:73  */
  assign n2384_o = n2371_o ? 1'b1 : n2383_o;
  assign n2385_o = n1909_o[84];
  /* TG68KdotC_Kernel.vhd:1731:73  */
  assign n2386_o = n2371_o ? 1'b1 : n2385_o;
  assign n2387_o = n1909_o[86];
  /* TG68KdotC_Kernel.vhd:1731:73  */
  assign n2388_o = n2371_o ? 1'b1 : n2387_o;
  /* TG68KdotC_Kernel.vhd:1731:73  */
  assign n2390_o = n2371_o ? 7'b0111110 : n2368_o;
  /* TG68KdotC_Kernel.vhd:1720:65  */
  assign n2391_o = n2355_o ? n2026_o : n2377_o;
  /* TG68KdotC_Kernel.vhd:1720:65  */
  assign n2393_o = n2355_o ? 1'b0 : n2380_o;
  assign n2394_o = n1909_o[26];
  /* TG68KdotC_Kernel.vhd:1720:65  */
  assign n2395_o = n2355_o ? n2394_o : n2382_o;
  assign n2396_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:1720:65  */
  assign n2397_o = n2355_o ? n2396_o : n2364_o;
  assign n2398_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:1720:65  */
  assign n2399_o = n2355_o ? n2398_o : n2384_o;
  /* TG68KdotC_Kernel.vhd:1720:65  */
  assign n2400_o = n2355_o ? n2358_o : n2366_o;
  assign n2401_o = n1909_o[84];
  /* TG68KdotC_Kernel.vhd:1720:65  */
  assign n2402_o = n2355_o ? n2401_o : n2386_o;
  assign n2403_o = n1909_o[86];
  /* TG68KdotC_Kernel.vhd:1720:65  */
  assign n2404_o = n2355_o ? n2403_o : n2388_o;
  /* TG68KdotC_Kernel.vhd:1720:65  */
  assign n2405_o = n2355_o ? n2360_o : n2390_o;
  /* TG68KdotC_Kernel.vhd:1712:57  */
  assign n2406_o = n2340_o ? n2350_o : n1921_o;
  /* TG68KdotC_Kernel.vhd:1712:57  */
  assign n2407_o = n2340_o ? n2391_o : n2026_o;
  /* TG68KdotC_Kernel.vhd:1712:57  */
  assign n2409_o = n2340_o ? n2393_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1712:57  */
  assign n2412_o = n2340_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1712:57  */
  assign n2415_o = n2340_o ? 1'b0 : 1'b1;
  assign n2416_o = n1909_o[26];
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2417_o = n2995_o ? n2395_o : n2416_o;
  assign n2418_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:1712:57  */
  assign n2419_o = n2340_o ? n2397_o : n2418_o;
  assign n2420_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2421_o = n2524_o ? n2399_o : n2420_o;
  assign n2422_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:1712:57  */
  assign n2423_o = n2340_o ? n2400_o : n2422_o;
  assign n2424_o = n1909_o[84];
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2425_o = n3017_o ? n2402_o : n2424_o;
  assign n2426_o = n1909_o[86];
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2427_o = n3019_o ? n2404_o : n2426_o;
  /* TG68KdotC_Kernel.vhd:1712:57  */
  assign n2428_o = n2340_o ? n2405_o : n2180_o;
  /* TG68KdotC_Kernel.vhd:1746:66  */
  assign n2429_o = opcode[10:9];
  /* TG68KdotC_Kernel.vhd:1746:79  */
  assign n2431_o = n2429_o != 2'b11;
  /* TG68KdotC_Kernel.vhd:1747:66  */
  assign n2432_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:1747:78  */
  assign n2434_o = n2432_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:1746:86  */
  assign n2435_o = n2434_o & n2431_o;
  /* TG68KdotC_Kernel.vhd:1747:95  */
  assign n2436_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1747:107  */
  assign n2438_o = n2436_o != 3'b011;
  /* TG68KdotC_Kernel.vhd:1747:85  */
  assign n2439_o = n2438_o & n2435_o;
  /* TG68KdotC_Kernel.vhd:1747:125  */
  assign n2440_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1747:137  */
  assign n2442_o = n2440_o != 3'b100;
  /* TG68KdotC_Kernel.vhd:1747:115  */
  assign n2443_o = n2442_o & n2439_o;
  /* TG68KdotC_Kernel.vhd:1747:155  */
  assign n2444_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:1747:167  */
  assign n2446_o = n2444_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:1747:145  */
  assign n2447_o = n2446_o & n2443_o;
  /* TG68KdotC_Kernel.vhd:1749:83  */
  assign n2449_o = opcode[10:9];
  assign n2452_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:1750:65  */
  assign n2453_o = decodeopc ? 1'b1 : n2452_o;
  assign n2454_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2455_o = n2500_o ? 1'b1 : n2454_o;
  /* TG68KdotC_Kernel.vhd:1750:65  */
  assign n2457_o = decodeopc ? 7'b0000001 : n2180_o;
  /* TG68KdotC_Kernel.vhd:1755:71  */
  assign n2458_o = set[62];
  assign n2461_o = n1909_o[39];
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2462_o = n2494_o ? 1'b1 : n2461_o;
  assign n2463_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2464_o = n2498_o ? 1'b1 : n2463_o;
  /* TG68KdotC_Kernel.vhd:1759:79  */
  assign n2466_o = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:1759:85  */
  assign n2467_o = nextpass & n2466_o;
  /* TG68KdotC_Kernel.vhd:1762:88  */
  assign n2470_o = exe_datatype != 2'b00;
  /* TG68KdotC_Kernel.vhd:1762:73  */
  assign n2473_o = n2470_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2475_o = n2483_o ? 2'b10 : n2026_o;
  /* TG68KdotC_Kernel.vhd:1759:65  */
  assign n2477_o = n2467_o ? n2473_o : 1'b0;
  assign n2478_o = n1909_o[82];
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2479_o = n2502_o ? 1'b1 : n2478_o;
  /* TG68KdotC_Kernel.vhd:1759:65  */
  assign n2481_o = n2467_o ? 7'b1001000 : n2457_o;
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2482_o = n2447_o ? n2449_o : n1921_o;
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2483_o = n2467_o & n2447_o;
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2486_o = n2447_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2489_o = n2447_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2491_o = n2447_o ? n2477_o : 1'b0;
  assign n2492_o = {1'b1, n2453_o};
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2494_o = n2458_o & n2447_o;
  assign n2495_o = n1909_o[43:42];
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2496_o = n2447_o ? n2492_o : n2495_o;
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2498_o = n2458_o & n2447_o;
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2500_o = decodeopc & n2447_o;
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2502_o = n2467_o & n2447_o;
  /* TG68KdotC_Kernel.vhd:1746:57  */
  assign n2503_o = n2447_o ? n2481_o : n2180_o;
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2504_o = n2319_o ? n2406_o : n2482_o;
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2505_o = n2319_o ? n2407_o : n2475_o;
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2507_o = n2319_o ? n2409_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2508_o = n2319_o ? n2412_o : n2486_o;
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2509_o = n2319_o ? n2415_o : n2489_o;
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2511_o = n2319_o ? 1'b0 : n2491_o;
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2513_o = n2340_o & n2319_o;
  assign n2514_o = n1909_o[39];
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2515_o = n2319_o ? n2514_o : n2462_o;
  assign n2516_o = n2496_o[0];
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2517_o = n2319_o ? n2419_o : n2516_o;
  assign n2518_o = n2496_o[1];
  assign n2519_o = n1909_o[43];
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2520_o = n2319_o ? n2519_o : n2518_o;
  assign n2521_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2522_o = n2319_o ? n2521_o : n2464_o;
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2524_o = n2340_o & n2319_o;
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2525_o = n2319_o ? n2423_o : n2455_o;
  assign n2526_o = n1909_o[82];
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2527_o = n2319_o ? n2526_o : n2479_o;
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2529_o = n2340_o & n2319_o;
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2531_o = n2340_o & n2319_o;
  /* TG68KdotC_Kernel.vhd:1711:49  */
  assign n2532_o = n2319_o ? n2428_o : n2503_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2533_o = n2979_o ? n2504_o : n1921_o;
  /* TG68KdotC_Kernel.vhd:1710:41  */
  assign n2534_o = n2318_o ? n2505_o : n2026_o;
  /* TG68KdotC_Kernel.vhd:1710:41  */
  assign n2536_o = n2318_o ? n2507_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1710:41  */
  assign n2538_o = n2318_o ? n2508_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1710:41  */
  assign n2540_o = n2318_o ? n2509_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1710:41  */
  assign n2542_o = n2318_o ? n2511_o : 1'b0;
  assign n2543_o = {n2520_o, n2517_o};
  assign n2544_o = {n2421_o, n2522_o};
  /* TG68KdotC_Kernel.vhd:1710:41  */
  assign n2546_o = n2513_o & n2318_o;
  assign n2547_o = n1909_o[39];
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2548_o = n2997_o ? n2515_o : n2547_o;
  assign n2549_o = n1909_o[43:42];
  /* TG68KdotC_Kernel.vhd:1710:41  */
  assign n2550_o = n2318_o ? n2543_o : n2549_o;
  assign n2551_o = n1909_o[56:55];
  /* TG68KdotC_Kernel.vhd:1710:41  */
  assign n2552_o = n2318_o ? n2544_o : n2551_o;
  assign n2553_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:1710:41  */
  assign n2554_o = n2318_o ? n2525_o : n2553_o;
  assign n2555_o = n1909_o[82];
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2556_o = n3015_o ? n2527_o : n2555_o;
  /* TG68KdotC_Kernel.vhd:1710:41  */
  assign n2558_o = n2529_o & n2318_o;
  /* TG68KdotC_Kernel.vhd:1710:41  */
  assign n2560_o = n2531_o & n2318_o;
  /* TG68KdotC_Kernel.vhd:1710:41  */
  assign n2561_o = n2318_o ? n2532_o : n2180_o;
  /* TG68KdotC_Kernel.vhd:1776:45  */
  assign n2562_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:1776:58  */
  assign n2564_o = n2562_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:1777:47  */
  assign n2565_o = cpu[0];
  /* TG68KdotC_Kernel.vhd:1777:65  */
  assign n2566_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:1777:77  */
  assign n2568_o = n2566_o != 2'b11;
  /* TG68KdotC_Kernel.vhd:1777:55  */
  assign n2569_o = n2568_o & n2565_o;
  /* TG68KdotC_Kernel.vhd:1777:94  */
  assign n2570_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:1777:106  */
  assign n2572_o = n2570_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:1777:84  */
  assign n2573_o = n2572_o & n2569_o;
  /* TG68KdotC_Kernel.vhd:1777:124  */
  assign n2574_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1777:136  */
  assign n2576_o = n2574_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:1777:153  */
  assign n2577_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:1777:165  */
  assign n2579_o = n2577_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1777:144  */
  assign n2580_o = n2576_o | n2579_o;
  /* TG68KdotC_Kernel.vhd:1777:113  */
  assign n2581_o = n2580_o & n2573_o;
  /* TG68KdotC_Kernel.vhd:1778:49  */
  assign n2584_o = svmode ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1778:49  */
  assign n2587_o = svmode ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1777:41  */
  assign n2589_o = n2581_o ? n2584_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1777:41  */
  assign n2591_o = n2581_o ? n2587_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1791:50  */
  assign n2592_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:1791:62  */
  assign n2594_o = n2592_o != 2'b11;
  /* TG68KdotC_Kernel.vhd:1791:79  */
  assign n2595_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1791:91  */
  assign n2597_o = n2595_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:1791:69  */
  assign n2598_o = n2597_o & n2594_o;
  /* TG68KdotC_Kernel.vhd:1792:58  */
  assign n2599_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:1792:71  */
  assign n2601_o = n2599_o == 3'b000;
  /* TG68KdotC_Kernel.vhd:1793:66  */
  assign n2602_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1793:78  */
  assign n2604_o = n2602_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:1793:95  */
  assign n2605_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:1793:107  */
  assign n2607_o = n2605_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1793:86  */
  assign n2608_o = n2604_o | n2607_o;
  /* TG68KdotC_Kernel.vhd:1793:123  */
  assign n2609_o = opcode[2:0];
  /* TG68KdotC_Kernel.vhd:1793:135  */
  assign n2611_o = n2609_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:1793:152  */
  assign n2612_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:1793:155  */
  assign n2613_o = ~n2612_o;
  /* TG68KdotC_Kernel.vhd:1793:142  */
  assign n2614_o = n2613_o & n2611_o;
  /* TG68KdotC_Kernel.vhd:1793:113  */
  assign n2615_o = n2608_o | n2614_o;
  /* TG68KdotC_Kernel.vhd:1793:57  */
  assign n2619_o = n2615_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1793:57  */
  assign n2622_o = n2615_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1793:57  */
  assign n2624_o = n2615_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1792:49  */
  assign n2626_o = n2601_o ? n2619_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1792:49  */
  assign n2628_o = n2601_o ? n2622_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1792:49  */
  assign n2630_o = n2601_o ? n2624_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1800:58  */
  assign n2631_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:1800:71  */
  assign n2633_o = n2631_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:1801:66  */
  assign n2634_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1801:78  */
  assign n2636_o = n2634_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:1801:95  */
  assign n2637_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:1801:107  */
  assign n2639_o = n2637_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1801:86  */
  assign n2640_o = n2636_o | n2639_o;
  /* TG68KdotC_Kernel.vhd:1801:123  */
  assign n2641_o = opcode[2:0];
  /* TG68KdotC_Kernel.vhd:1801:135  */
  assign n2643_o = n2641_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:1801:152  */
  assign n2644_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:1801:155  */
  assign n2645_o = ~n2644_o;
  /* TG68KdotC_Kernel.vhd:1801:142  */
  assign n2646_o = n2645_o & n2643_o;
  /* TG68KdotC_Kernel.vhd:1801:113  */
  assign n2647_o = n2640_o | n2646_o;
  /* TG68KdotC_Kernel.vhd:1801:57  */
  assign n2650_o = n2647_o ? n2626_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1801:57  */
  assign n2652_o = n2647_o ? n2628_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1801:57  */
  assign n2654_o = n2647_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1800:49  */
  assign n2655_o = n2633_o ? n2650_o : n2626_o;
  /* TG68KdotC_Kernel.vhd:1800:49  */
  assign n2656_o = n2633_o ? n2652_o : n2628_o;
  /* TG68KdotC_Kernel.vhd:1800:49  */
  assign n2658_o = n2633_o ? n2654_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1808:58  */
  assign n2659_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:1808:71  */
  assign n2661_o = n2659_o == 3'b010;
  /* TG68KdotC_Kernel.vhd:1808:87  */
  assign n2662_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:1808:100  */
  assign n2664_o = n2662_o == 3'b011;
  /* TG68KdotC_Kernel.vhd:1808:78  */
  assign n2665_o = n2661_o | n2664_o;
  /* TG68KdotC_Kernel.vhd:1809:66  */
  assign n2666_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1809:78  */
  assign n2668_o = n2666_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:1809:95  */
  assign n2669_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:1809:107  */
  assign n2671_o = n2669_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1809:86  */
  assign n2672_o = n2668_o | n2671_o;
  /* TG68KdotC_Kernel.vhd:1809:57  */
  assign n2675_o = n2672_o ? n2655_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1809:57  */
  assign n2677_o = n2672_o ? n2656_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1809:57  */
  assign n2679_o = n2672_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1808:49  */
  assign n2680_o = n2665_o ? n2675_o : n2655_o;
  /* TG68KdotC_Kernel.vhd:1808:49  */
  assign n2681_o = n2665_o ? n2677_o : n2656_o;
  /* TG68KdotC_Kernel.vhd:1808:49  */
  assign n2683_o = n2665_o ? n2679_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1816:58  */
  assign n2684_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:1816:71  */
  assign n2686_o = n2684_o == 3'b101;
  /* TG68KdotC_Kernel.vhd:1817:66  */
  assign n2687_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1817:78  */
  assign n2689_o = n2687_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:1817:95  */
  assign n2690_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:1817:107  */
  assign n2692_o = n2690_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1817:86  */
  assign n2693_o = n2689_o | n2692_o;
  /* TG68KdotC_Kernel.vhd:1817:123  */
  assign n2694_o = opcode[2:0];
  /* TG68KdotC_Kernel.vhd:1817:135  */
  assign n2696_o = n2694_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:1817:152  */
  assign n2697_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:1817:155  */
  assign n2698_o = ~n2697_o;
  /* TG68KdotC_Kernel.vhd:1817:142  */
  assign n2699_o = n2698_o & n2696_o;
  /* TG68KdotC_Kernel.vhd:1817:113  */
  assign n2700_o = n2693_o | n2699_o;
  /* TG68KdotC_Kernel.vhd:1817:57  */
  assign n2703_o = n2700_o ? n2680_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1817:57  */
  assign n2705_o = n2700_o ? n2681_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1817:57  */
  assign n2707_o = n2700_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1816:49  */
  assign n2708_o = n2686_o ? n2703_o : n2680_o;
  /* TG68KdotC_Kernel.vhd:1816:49  */
  assign n2709_o = n2686_o ? n2705_o : n2681_o;
  /* TG68KdotC_Kernel.vhd:1816:49  */
  assign n2711_o = n2686_o ? n2707_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1824:58  */
  assign n2712_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:1824:71  */
  assign n2714_o = n2712_o == 3'b110;
  /* TG68KdotC_Kernel.vhd:1825:66  */
  assign n2715_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1825:78  */
  assign n2717_o = n2715_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:1825:95  */
  assign n2718_o = opcode[2];
  /* TG68KdotC_Kernel.vhd:1825:98  */
  assign n2719_o = ~n2718_o;
  /* TG68KdotC_Kernel.vhd:1825:86  */
  assign n2720_o = n2717_o | n2719_o;
  /* TG68KdotC_Kernel.vhd:1825:57  */
  assign n2723_o = n2720_o ? n2708_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1825:57  */
  assign n2725_o = n2720_o ? n2709_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1825:57  */
  assign n2727_o = n2720_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1824:49  */
  assign n2728_o = n2714_o ? n2723_o : n2708_o;
  /* TG68KdotC_Kernel.vhd:1824:49  */
  assign n2729_o = n2714_o ? n2725_o : n2709_o;
  /* TG68KdotC_Kernel.vhd:1824:49  */
  assign n2731_o = n2714_o ? n2727_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1832:61  */
  assign n2732_o = set_exec[5];
  /* TG68KdotC_Kernel.vhd:1832:80  */
  assign n2733_o = set_exec[6];
  /* TG68KdotC_Kernel.vhd:1832:69  */
  assign n2734_o = n2732_o | n2733_o;
  /* TG68KdotC_Kernel.vhd:1832:100  */
  assign n2735_o = set_exec[3];
  /* TG68KdotC_Kernel.vhd:1832:89  */
  assign n2736_o = n2734_o | n2735_o;
  /* TG68KdotC_Kernel.vhd:1832:120  */
  assign n2737_o = set_exec[7];
  /* TG68KdotC_Kernel.vhd:1832:109  */
  assign n2738_o = n2736_o | n2737_o;
  /* TG68KdotC_Kernel.vhd:1832:140  */
  assign n2739_o = set_exec[8];
  /* TG68KdotC_Kernel.vhd:1832:129  */
  assign n2740_o = n2738_o | n2739_o;
  /* TG68KdotC_Kernel.vhd:1833:66  */
  assign n2741_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:1833:69  */
  assign n2742_o = ~n2741_o;
  /* TG68KdotC_Kernel.vhd:1833:84  */
  assign n2743_o = opcode[5:0];
  /* TG68KdotC_Kernel.vhd:1833:96  */
  assign n2745_o = n2743_o == 6'b111100;
  /* TG68KdotC_Kernel.vhd:1833:74  */
  assign n2746_o = n2745_o & n2742_o;
  /* TG68KdotC_Kernel.vhd:1833:119  */
  assign n2747_o = set_exec[6];
  /* TG68KdotC_Kernel.vhd:1833:139  */
  assign n2748_o = set_exec[5];
  /* TG68KdotC_Kernel.vhd:1833:128  */
  assign n2749_o = n2747_o | n2748_o;
  /* TG68KdotC_Kernel.vhd:1833:158  */
  assign n2750_o = set_exec[7];
  /* TG68KdotC_Kernel.vhd:1833:147  */
  assign n2751_o = n2749_o | n2750_o;
  /* TG68KdotC_Kernel.vhd:1833:106  */
  assign n2752_o = n2751_o & n2746_o;
  /* TG68KdotC_Kernel.vhd:1834:92  */
  assign n2753_o = ~svmode;
  /* TG68KdotC_Kernel.vhd:1834:82  */
  assign n2754_o = n2753_o & decodeopc;
  /* TG68KdotC_Kernel.vhd:1834:107  */
  assign n2755_o = opcode[6];
  /* TG68KdotC_Kernel.vhd:1834:97  */
  assign n2756_o = n2755_o & n2754_o;
  /* TG68KdotC_Kernel.vhd:1840:90  */
  assign n2758_o = opcode[6];
  assign n2760_o = n1909_o[52];
  /* TG68KdotC_Kernel.vhd:1840:81  */
  assign n2761_o = n2758_o ? 1'b1 : n2760_o;
  /* TG68KdotC_Kernel.vhd:1844:104  */
  assign n2763_o = set_exec[6];
  /* TG68KdotC_Kernel.vhd:1845:104  */
  assign n2764_o = set_exec[7];
  /* TG68KdotC_Kernel.vhd:1846:103  */
  assign n2765_o = set_exec[5];
  /* TG68KdotC_Kernel.vhd:1839:73  */
  assign n2767_o = decodeopc ? 2'b01 : n2026_o;
  assign n2768_o = {n2765_o, n2764_o, n2763_o};
  assign n2769_o = {n2761_o, 1'b1};
  assign n2770_o = n1909_o[19:17];
  /* TG68KdotC_Kernel.vhd:1839:73  */
  assign n2771_o = decodeopc ? n2768_o : n2770_o;
  assign n2772_o = n1909_o[52:51];
  /* TG68KdotC_Kernel.vhd:1839:73  */
  assign n2773_o = decodeopc ? n2769_o : n2772_o;
  /* TG68KdotC_Kernel.vhd:1839:73  */
  assign n2775_o = decodeopc ? 7'b0011000 : n2180_o;
  /* TG68KdotC_Kernel.vhd:1834:65  */
  assign n2776_o = n2756_o ? n2026_o : n2767_o;
  /* TG68KdotC_Kernel.vhd:1834:65  */
  assign n2779_o = n2756_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1834:65  */
  assign n2781_o = n2756_o ? 1'b1 : n2729_o;
  assign n2782_o = n1909_o[19:17];
  /* TG68KdotC_Kernel.vhd:1834:65  */
  assign n2783_o = n2756_o ? n2782_o : n2771_o;
  assign n2784_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:1834:65  */
  assign n2785_o = n2756_o ? n2784_o : 1'b1;
  assign n2786_o = n1909_o[52:51];
  /* TG68KdotC_Kernel.vhd:1834:65  */
  assign n2787_o = n2756_o ? n2786_o : n2773_o;
  /* TG68KdotC_Kernel.vhd:1834:65  */
  assign n2788_o = n2756_o ? n2180_o : n2775_o;
  /* TG68KdotC_Kernel.vhd:1851:69  */
  assign n2789_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:1851:72  */
  assign n2790_o = ~n2789_o;
  /* TG68KdotC_Kernel.vhd:1851:86  */
  assign n2791_o = opcode[5:0];
  /* TG68KdotC_Kernel.vhd:1851:98  */
  assign n2793_o = n2791_o != 6'b111100;
  /* TG68KdotC_Kernel.vhd:1851:77  */
  assign n2794_o = n2790_o | n2793_o;
  /* TG68KdotC_Kernel.vhd:1851:121  */
  assign n2795_o = set_exec[6];
  /* TG68KdotC_Kernel.vhd:1851:141  */
  assign n2796_o = set_exec[5];
  /* TG68KdotC_Kernel.vhd:1851:130  */
  assign n2797_o = n2795_o | n2796_o;
  /* TG68KdotC_Kernel.vhd:1851:160  */
  assign n2798_o = set_exec[7];
  /* TG68KdotC_Kernel.vhd:1851:149  */
  assign n2799_o = n2797_o | n2798_o;
  /* TG68KdotC_Kernel.vhd:1851:169  */
  assign n2800_o = ~n2799_o;
  /* TG68KdotC_Kernel.vhd:1851:109  */
  assign n2801_o = n2794_o | n2800_o;
  /* TG68KdotC_Kernel.vhd:1857:84  */
  assign n2805_o = datatype == 2'b10;
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2807_o = n2856_o ? 1'b1 : n2171_o;
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2809_o = n2845_o ? 1'b1 : n2154_o;
  assign n2810_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2811_o = n2851_o ? 1'b1 : n2810_o;
  assign n2812_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2813_o = n2855_o ? 1'b1 : n2812_o;
  /* TG68KdotC_Kernel.vhd:1852:65  */
  assign n2814_o = n2805_o & decodeopc;
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2816_o = n2861_o ? 7'b0011101 : n2180_o;
  /* TG68KdotC_Kernel.vhd:1861:74  */
  assign n2817_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:1861:86  */
  assign n2819_o = n2817_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:1861:65  */
  assign n2822_o = n2819_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1864:74  */
  assign n2823_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:1864:87  */
  assign n2825_o = n2823_o != 3'b110;
  /* TG68KdotC_Kernel.vhd:1865:82  */
  assign n2826_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:1865:94  */
  assign n2828_o = n2826_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1865:73  */
  assign n2831_o = n2828_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1864:65  */
  assign n2834_o = n2825_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1864:65  */
  assign n2836_o = n2825_o ? n2831_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1870:74  */
  assign n2837_o = opcode[10:9];
  /* TG68KdotC_Kernel.vhd:1870:87  */
  assign n2839_o = n2837_o == 2'b10;
  assign n2841_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2842_o = n2853_o ? 1'b1 : n2841_o;
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2844_o = n2801_o ? n2834_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2845_o = decodeopc & n2801_o;
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2847_o = n2801_o ? n2728_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2849_o = n2801_o ? n2729_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2851_o = decodeopc & n2801_o;
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2853_o = n2839_o & n2801_o;
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2855_o = decodeopc & n2801_o;
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2856_o = n2814_o & n2801_o;
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2858_o = n2801_o ? n2822_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2860_o = n2801_o ? n2836_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1851:57  */
  assign n2861_o = decodeopc & n2801_o;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2862_o = n2916_o ? n2776_o : n2026_o;
  /* TG68KdotC_Kernel.vhd:1833:57  */
  assign n2864_o = n2752_o ? 1'b0 : n2844_o;
  /* TG68KdotC_Kernel.vhd:1833:57  */
  assign n2865_o = n2752_o ? n2154_o : n2809_o;
  /* TG68KdotC_Kernel.vhd:1833:57  */
  assign n2866_o = n2752_o ? n2728_o : n2847_o;
  /* TG68KdotC_Kernel.vhd:1833:57  */
  assign n2868_o = n2752_o ? n2779_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1833:57  */
  assign n2869_o = n2752_o ? n2781_o : n2849_o;
  assign n2870_o = n1909_o[19:17];
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2871_o = n2927_o ? n2783_o : n2870_o;
  assign n2872_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:1833:57  */
  assign n2873_o = n2752_o ? n2872_o : n2811_o;
  assign n2874_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2875_o = n2931_o ? n2785_o : n2874_o;
  assign n2876_o = n1909_o[52:51];
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2877_o = n2933_o ? n2787_o : n2876_o;
  assign n2878_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:1833:57  */
  assign n2879_o = n2752_o ? n2878_o : n2842_o;
  assign n2880_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:1833:57  */
  assign n2881_o = n2752_o ? n2880_o : n2813_o;
  /* TG68KdotC_Kernel.vhd:1833:57  */
  assign n2882_o = n2752_o ? n2171_o : n2807_o;
  /* TG68KdotC_Kernel.vhd:1833:57  */
  assign n2884_o = n2752_o ? 1'b0 : n2858_o;
  /* TG68KdotC_Kernel.vhd:1833:57  */
  assign n2886_o = n2752_o ? 1'b0 : n2860_o;
  /* TG68KdotC_Kernel.vhd:1833:57  */
  assign n2887_o = n2752_o ? n2788_o : n2816_o;
  /* TG68KdotC_Kernel.vhd:1832:49  */
  assign n2888_o = n2752_o & n2740_o;
  /* TG68KdotC_Kernel.vhd:1832:49  */
  assign n2890_o = n2740_o ? n2864_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2891_o = n2919_o ? n2865_o : n2154_o;
  /* TG68KdotC_Kernel.vhd:1832:49  */
  assign n2893_o = n2740_o ? n2866_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1832:49  */
  assign n2895_o = n2740_o ? n2868_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1832:49  */
  assign n2897_o = n2740_o ? n2869_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1832:49  */
  assign n2899_o = n2752_o & n2740_o;
  assign n2900_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2901_o = n2929_o ? n2873_o : n2900_o;
  /* TG68KdotC_Kernel.vhd:1832:49  */
  assign n2903_o = n2752_o & n2740_o;
  /* TG68KdotC_Kernel.vhd:1832:49  */
  assign n2905_o = n2752_o & n2740_o;
  assign n2906_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2907_o = n2935_o ? n2879_o : n2906_o;
  assign n2908_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2909_o = n2937_o ? n2881_o : n2908_o;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2910_o = n2938_o ? n2882_o : n2171_o;
  /* TG68KdotC_Kernel.vhd:1832:49  */
  assign n2912_o = n2740_o ? n2884_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1832:49  */
  assign n2914_o = n2740_o ? n2886_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2915_o = n2948_o ? n2887_o : n2180_o;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2916_o = n2888_o & n2598_o;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2918_o = n2598_o ? n2890_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2919_o = n2740_o & n2598_o;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2921_o = n2598_o ? n2893_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2923_o = n2598_o ? n2895_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2925_o = n2598_o ? n2897_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2927_o = n2899_o & n2598_o;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2929_o = n2740_o & n2598_o;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2931_o = n2903_o & n2598_o;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2933_o = n2905_o & n2598_o;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2935_o = n2740_o & n2598_o;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2937_o = n2740_o & n2598_o;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2938_o = n2740_o & n2598_o;
  assign n2939_o = {n2731_o, n2711_o, n2658_o, n2630_o};
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2941_o = n2598_o ? n2683_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2943_o = n2598_o ? n2939_o : 4'b0000;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2945_o = n2598_o ? n2912_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2947_o = n2598_o ? n2914_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1791:41  */
  assign n2948_o = n2740_o & n2598_o;
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2949_o = n2564_o ? n2026_o : n2862_o;
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2951_o = n2564_o ? 1'b0 : n2918_o;
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2952_o = n2564_o ? n2154_o : n2891_o;
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2953_o = n2564_o ? n2589_o : n2921_o;
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2954_o = n2564_o ? n2591_o : n2923_o;
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2956_o = n2564_o ? 1'b1 : n2925_o;
  assign n2957_o = n1909_o[19:17];
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2958_o = n2564_o ? n2957_o : n2871_o;
  assign n2959_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2960_o = n2564_o ? n2959_o : n2901_o;
  assign n2961_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2962_o = n2564_o ? n2961_o : n2875_o;
  assign n2963_o = n1909_o[52:51];
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2964_o = n2564_o ? n2963_o : n2877_o;
  assign n2965_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2966_o = n2564_o ? n2965_o : n2907_o;
  assign n2967_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2968_o = n2564_o ? n2967_o : n2909_o;
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2969_o = n2564_o ? n2171_o : n2910_o;
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2971_o = n2564_o ? 1'b0 : n2941_o;
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2973_o = n2564_o ? 4'b0000 : n2943_o;
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2975_o = n2564_o ? 1'b0 : n2945_o;
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2977_o = n2564_o ? 1'b0 : n2947_o;
  /* TG68KdotC_Kernel.vhd:1776:33  */
  assign n2978_o = n2564_o ? n2180_o : n2915_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2979_o = n2318_o & n2317_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2980_o = n2317_o ? n2534_o : n2949_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2982_o = n2317_o ? 1'b0 : n2951_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2984_o = n2317_o ? n2536_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2985_o = n2317_o ? n2154_o : n2952_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2986_o = n2317_o ? n2538_o : n2953_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2988_o = n2317_o ? 1'b0 : n2954_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2989_o = n2317_o ? n2540_o : n2956_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2991_o = n2317_o ? n2542_o : 1'b0;
  assign n2992_o = n1909_o[19:17];
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2993_o = n2317_o ? n2992_o : n2958_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2995_o = n2546_o & n2317_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2997_o = n2318_o & n2317_o;
  assign n2998_o = n2550_o[0];
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n2999_o = n2317_o ? n2998_o : n2960_o;
  assign n3000_o = n2550_o[1];
  assign n3001_o = n1909_o[43];
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3002_o = n2317_o ? n3000_o : n3001_o;
  assign n3003_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3004_o = n2317_o ? n3003_o : n2962_o;
  assign n3005_o = n1909_o[52:51];
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3006_o = n2317_o ? n3005_o : n2964_o;
  assign n3007_o = n2552_o[0];
  assign n3008_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3009_o = n2317_o ? n3007_o : n3008_o;
  assign n3010_o = n2552_o[1];
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3011_o = n2317_o ? n3010_o : n2966_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3012_o = n2317_o ? n2554_o : n2968_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3013_o = n2317_o ? n2171_o : n2969_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3015_o = n2318_o & n2317_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3017_o = n2558_o & n2317_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3019_o = n2560_o & n2317_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3021_o = n2317_o ? 1'b0 : n2971_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3023_o = n2317_o ? 4'b0000 : n2973_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3025_o = n2317_o ? 1'b0 : n2975_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3027_o = n2317_o ? 1'b0 : n2977_o;
  /* TG68KdotC_Kernel.vhd:1709:33  */
  assign n3028_o = n2317_o ? n2561_o : n2978_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3029_o = n2222_o ? n2293_o : n2533_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3030_o = n2222_o ? n2026_o : n2980_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3031_o = n2222_o ? n2295_o : n2982_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3033_o = n2222_o ? 1'b0 : n2984_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3034_o = n2222_o ? n2154_o : n2985_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3035_o = n2222_o ? n2298_o : n2986_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3037_o = n2222_o ? 1'b0 : n2988_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3038_o = n2222_o ? n2301_o : n2989_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3040_o = n2222_o ? n2303_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3042_o = n2222_o ? 1'b0 : n2991_o;
  assign n3043_o = {n3002_o, n2999_o};
  assign n3044_o = {n3011_o, n3009_o};
  assign n3045_o = n1909_o[19:17];
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3046_o = n2222_o ? n3045_o : n2993_o;
  assign n3047_o = n1909_o[26];
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3048_o = n2222_o ? n3047_o : n2417_o;
  assign n3049_o = n1909_o[39];
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3050_o = n2222_o ? n3049_o : n2548_o;
  assign n3051_o = n3043_o[0];
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3052_o = n2222_o ? n2280_o : n3051_o;
  assign n3053_o = n3043_o[1];
  assign n3054_o = n1909_o[43];
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3055_o = n2222_o ? n3054_o : n3053_o;
  assign n3056_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3057_o = n2222_o ? n3056_o : n3004_o;
  assign n3058_o = n1909_o[52:51];
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3059_o = n2222_o ? n3058_o : n3006_o;
  assign n3060_o = n1909_o[56:55];
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3061_o = n2222_o ? n3060_o : n3044_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3062_o = n2222_o ? n2282_o : n3012_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3063_o = n2222_o ? n2171_o : n3013_o;
  assign n3064_o = n1909_o[82];
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3065_o = n2222_o ? n3064_o : n2556_o;
  assign n3066_o = n1909_o[84];
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3067_o = n2222_o ? n3066_o : n2425_o;
  assign n3068_o = n1909_o[86];
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3069_o = n2222_o ? n3068_o : n2427_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3071_o = n2222_o ? 1'b0 : n3021_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3073_o = n2222_o ? 4'b0000 : n3023_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3075_o = n2222_o ? n2309_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3076_o = n2222_o ? n2311_o : n3025_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3077_o = n2222_o ? n2313_o : n3027_o;
  /* TG68KdotC_Kernel.vhd:1678:33  */
  assign n3078_o = n2222_o ? n2284_o : n3028_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3080_o = n2190_o ? 2'b00 : n3029_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3081_o = n2190_o ? n2026_o : n3030_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3083_o = n2190_o ? 1'b0 : n3031_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3085_o = n2190_o ? 1'b0 : n3033_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3087_o = n2190_o ? n2217_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3088_o = n2190_o ? n2210_o : n3034_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3090_o = n2190_o ? 1'b0 : n3035_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3092_o = n2190_o ? 1'b0 : n3037_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3094_o = n2190_o ? 1'b0 : n3038_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3096_o = n2190_o ? 1'b0 : n3040_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3098_o = n2190_o ? 1'b0 : n3042_o;
  assign n3099_o = {n3055_o, n3052_o};
  assign n3100_o = {1'b1, 1'b1};
  assign n3101_o = n1909_o[19:17];
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3102_o = n2190_o ? n3101_o : n3046_o;
  assign n3103_o = n1909_o[26];
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3104_o = n2190_o ? n3103_o : n3048_o;
  assign n3105_o = n1909_o[37];
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3106_o = n2190_o ? n2206_o : n3105_o;
  assign n3107_o = n1909_o[39];
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3108_o = n2190_o ? n3107_o : n3050_o;
  assign n3109_o = n1909_o[43:42];
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3110_o = n2190_o ? n3109_o : n3099_o;
  assign n3111_o = n3100_o[0];
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3112_o = n2190_o ? n3111_o : n3057_o;
  assign n3113_o = n3100_o[1];
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3114_o = n2190_o ? n3113_o : n2168_o;
  assign n3115_o = n1909_o[52:51];
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3116_o = n2190_o ? n3115_o : n3059_o;
  assign n3117_o = n1909_o[56:55];
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3118_o = n2190_o ? n3117_o : n3061_o;
  assign n3119_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3120_o = n2190_o ? n3119_o : n3062_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3121_o = n2190_o ? n2171_o : n3063_o;
  assign n3122_o = n1909_o[82];
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3123_o = n2190_o ? n3122_o : n3065_o;
  assign n3124_o = n1909_o[84];
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3125_o = n2190_o ? n3124_o : n3067_o;
  assign n3126_o = n1909_o[86];
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3127_o = n2190_o ? n3126_o : n3069_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3129_o = n2190_o ? n2201_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3131_o = n2190_o ? 1'b0 : n3071_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3133_o = n2190_o ? 4'b0000 : n3073_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3135_o = n2190_o ? 1'b0 : n3075_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3137_o = n2190_o ? 1'b0 : n3076_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3138_o = n2190_o ? n2203_o : n3077_o;
  /* TG68KdotC_Kernel.vhd:1656:25  */
  assign n3139_o = n2190_o ? n2214_o : n3078_o;
  /* TG68KdotC_Kernel.vhd:1655:25  */
  assign n3141_o = n2185_o == 4'b0000;
  /* TG68KdotC_Kernel.vhd:1890:44  */
  assign n3142_o = opcode[11:10];
  /* TG68KdotC_Kernel.vhd:1890:58  */
  assign n3144_o = n3142_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1890:73  */
  assign n3145_o = opcode[8:6];
  /* TG68KdotC_Kernel.vhd:1890:85  */
  assign n3147_o = n3145_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:1890:64  */
  assign n3148_o = n3144_o | n3147_o;
  /* TG68KdotC_Kernel.vhd:1891:43  */
  assign n3149_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:1891:55  */
  assign n3151_o = n3149_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:1891:73  */
  assign n3152_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:1891:85  */
  assign n3154_o = n3152_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1891:64  */
  assign n3155_o = n3151_o | n3154_o;
  /* TG68KdotC_Kernel.vhd:1890:94  */
  assign n3156_o = n3155_o & n3148_o;
  /* TG68KdotC_Kernel.vhd:1892:43  */
  assign n3157_o = opcode[13];
  /* TG68KdotC_Kernel.vhd:1892:62  */
  assign n3158_o = opcode[8:6];
  /* TG68KdotC_Kernel.vhd:1892:74  */
  assign n3160_o = n3158_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:1892:92  */
  assign n3161_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1892:104  */
  assign n3163_o = n3161_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:1892:82  */
  assign n3164_o = n3163_o & n3160_o;
  /* TG68KdotC_Kernel.vhd:1892:52  */
  assign n3165_o = n3157_o | n3164_o;
  /* TG68KdotC_Kernel.vhd:1891:92  */
  assign n3166_o = n3165_o & n3156_o;
  /* TG68KdotC_Kernel.vhd:1895:50  */
  assign n3168_o = opcode[8:6];
  /* TG68KdotC_Kernel.vhd:1895:62  */
  assign n3170_o = n3168_o == 3'b001;
  assign n3172_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:1895:41  */
  assign n3173_o = n3170_o ? 1'b1 : n3172_o;
  /* TG68KdotC_Kernel.vhd:1898:50  */
  assign n3174_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:1898:62  */
  assign n3176_o = n3174_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1899:58  */
  assign n3177_o = opcode[8:7];
  /* TG68KdotC_Kernel.vhd:1899:70  */
  assign n3179_o = n3177_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1899:49  */
  assign n3182_o = n3179_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1898:41  */
  assign n3184_o = n3176_o ? n3182_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1903:52  */
  assign n3185_o = opcode[13:12];
  /* TG68KdotC_Kernel.vhd:1904:49  */
  assign n3187_o = n3185_o == 2'b01;
  /* TG68KdotC_Kernel.vhd:1905:49  */
  assign n3189_o = n3185_o == 2'b10;
  assign n3190_o = {n3189_o, n3187_o};
  /* TG68KdotC_Kernel.vhd:1903:41  */
  always @*
    case (n3190_o)
      2'b10: n3194_o = 2'b10;
      2'b01: n3194_o = 2'b00;
      default: n3194_o = 2'b01;
    endcase
  /* TG68KdotC_Kernel.vhd:1909:50  */
  assign n3195_o = opcode[3];
  /* TG68KdotC_Kernel.vhd:1909:41  */
  assign n3198_o = n3195_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1913:66  */
  assign n3199_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:1913:78  */
  assign n3201_o = n3199_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1913:57  */
  assign n3202_o = nextpass | n3201_o;
  /* TG68KdotC_Kernel.vhd:1915:58  */
  assign n3203_o = opcode[8:6];
  /* TG68KdotC_Kernel.vhd:1915:70  */
  assign n3205_o = n3203_o != 3'b000;
  /* TG68KdotC_Kernel.vhd:1915:49  */
  assign n3208_o = n3205_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1913:41  */
  assign n3210_o = n3202_o ? n3208_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1913:41  */
  assign n3213_o = n3202_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1920:55  */
  assign n3215_o = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:1920:89  */
  assign n3216_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:1920:101  */
  assign n3218_o = n3216_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:1920:107  */
  assign n3219_o = decodeopc & n3218_o;
  /* TG68KdotC_Kernel.vhd:1920:79  */
  assign n3220_o = nextpass | n3219_o;
  /* TG68KdotC_Kernel.vhd:1920:61  */
  assign n3221_o = n3220_o & n3215_o;
  /* TG68KdotC_Kernel.vhd:1921:60  */
  assign n3222_o = opcode[8:6];
  /* TG68KdotC_Kernel.vhd:1922:57  */
  assign n3225_o = n3222_o == 3'b000;
  /* TG68KdotC_Kernel.vhd:1922:67  */
  assign n3227_o = n3222_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:1922:67  */
  assign n3228_o = n3225_o | n3227_o;
  /* TG68KdotC_Kernel.vhd:1925:74  */
  assign n3229_o = opcode[6];
  /* TG68KdotC_Kernel.vhd:1927:82  */
  assign n3231_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:1927:95  */
  assign n3233_o = n3231_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:1925:65  */
  assign n3235_o = n3240_o ? 1'b1 : n2168_o;
  assign n3236_o = n2162_o[0];
  assign n3237_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n3238_o = n2037_o ? n3236_o : n3237_o;
  /* TG68KdotC_Kernel.vhd:1925:65  */
  assign n3239_o = n3229_o ? 1'b1 : n3238_o;
  /* TG68KdotC_Kernel.vhd:1925:65  */
  assign n3240_o = n3233_o & n3229_o;
  /* TG68KdotC_Kernel.vhd:1931:74  */
  assign n3241_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:1933:82  */
  assign n3243_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:1933:95  */
  assign n3245_o = n3243_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:1931:65  */
  assign n3247_o = n3252_o ? 1'b1 : n3235_o;
  assign n3248_o = n2162_o[1];
  assign n3249_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n3250_o = n2037_o ? n3248_o : n3249_o;
  /* TG68KdotC_Kernel.vhd:1931:65  */
  assign n3251_o = n3241_o ? 1'b1 : n3250_o;
  /* TG68KdotC_Kernel.vhd:1931:65  */
  assign n3252_o = n3245_o & n3241_o;
  /* TG68KdotC_Kernel.vhd:1939:76  */
  assign n3253_o = ~nextpass;
  assign n3255_o = n1909_o[40];
  /* TG68KdotC_Kernel.vhd:1939:65  */
  assign n3256_o = n3253_o ? 1'b1 : n3255_o;
  /* TG68KdotC_Kernel.vhd:1924:57  */
  assign n3258_o = n3222_o == 3'b010;
  /* TG68KdotC_Kernel.vhd:1924:67  */
  assign n3260_o = n3222_o == 3'b011;
  /* TG68KdotC_Kernel.vhd:1924:67  */
  assign n3261_o = n3258_o | n3260_o;
  /* TG68KdotC_Kernel.vhd:1924:73  */
  assign n3263_o = n3222_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:1924:73  */
  assign n3264_o = n3261_o | n3263_o;
  /* TG68KdotC_Kernel.vhd:1942:57  */
  assign n3266_o = n3222_o == 3'b101;
  /* TG68KdotC_Kernel.vhd:1945:57  */
  assign n3268_o = n3222_o == 3'b110;
  /* TG68KdotC_Kernel.vhd:1949:76  */
  assign n3269_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:1950:73  */
  assign n3271_o = n3269_o == 3'b000;
  /* TG68KdotC_Kernel.vhd:1952:73  */
  assign n3274_o = n3269_o == 3'b001;
  assign n3275_o = {n3274_o, n3271_o};
  /* TG68KdotC_Kernel.vhd:1949:65  */
  always @*
    case (n3275_o)
      2'b10: n3276_o = 1'b1;
      2'b01: n3276_o = n2171_o;
      default: n3276_o = n2171_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1949:65  */
  always @*
    case (n3275_o)
      2'b10: n3279_o = 7'b0000011;
      2'b01: n3279_o = 7'b0000011;
      default: n3279_o = n2180_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1948:57  */
  assign n3281_o = n3222_o == 3'b111;
  assign n3282_o = {n3281_o, n3268_o, n3266_o, n3264_o, n3228_o};
  /* TG68KdotC_Kernel.vhd:1921:49  */
  always @*
    case (n3282_o)
      5'b10000: n3284_o = n2026_o;
      5'b01000: n3284_o = n2026_o;
      5'b00100: n3284_o = n2026_o;
      5'b00010: n3284_o = 2'b11;
      5'b00001: n3284_o = n2026_o;
      default: n3284_o = n2026_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1921:49  */
  always @*
    case (n3282_o)
      5'b10000: n3286_o = n2151_o;
      5'b01000: n3286_o = 1'b1;
      5'b00100: n3286_o = n2151_o;
      5'b00010: n3286_o = n2151_o;
      5'b00001: n3286_o = n2151_o;
      default: n3286_o = n2151_o;
    endcase
  assign n3287_o = n1909_o[40];
  /* TG68KdotC_Kernel.vhd:1921:49  */
  always @*
    case (n3282_o)
      5'b10000: n3288_o = n3287_o;
      5'b01000: n3288_o = n3287_o;
      5'b00100: n3288_o = n3287_o;
      5'b00010: n3288_o = n3256_o;
      5'b00001: n3288_o = n3287_o;
      default: n3288_o = n3287_o;
    endcase
  assign n3289_o = n2162_o[0];
  assign n3290_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n3291_o = n2037_o ? n3289_o : n3290_o;
  /* TG68KdotC_Kernel.vhd:1921:49  */
  always @*
    case (n3282_o)
      5'b10000: n3292_o = n3291_o;
      5'b01000: n3292_o = n3291_o;
      5'b00100: n3292_o = n3291_o;
      5'b00010: n3292_o = n3239_o;
      5'b00001: n3292_o = n3291_o;
      default: n3292_o = n3291_o;
    endcase
  assign n3293_o = n2162_o[1];
  assign n3294_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n3295_o = n2037_o ? n3293_o : n3294_o;
  /* TG68KdotC_Kernel.vhd:1921:49  */
  always @*
    case (n3282_o)
      5'b10000: n3296_o = n3295_o;
      5'b01000: n3296_o = n3295_o;
      5'b00100: n3296_o = n3295_o;
      5'b00010: n3296_o = n3251_o;
      5'b00001: n3296_o = n3295_o;
      default: n3296_o = n3295_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1921:49  */
  always @*
    case (n3282_o)
      5'b10000: n3297_o = n2168_o;
      5'b01000: n3297_o = n2168_o;
      5'b00100: n3297_o = n2168_o;
      5'b00010: n3297_o = n3247_o;
      5'b00001: n3297_o = n2168_o;
      default: n3297_o = n2168_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1921:49  */
  always @*
    case (n3282_o)
      5'b10000: n3298_o = n3276_o;
      5'b01000: n3298_o = n2171_o;
      5'b00100: n3298_o = n2171_o;
      5'b00010: n3298_o = n2171_o;
      5'b00001: n3298_o = n2171_o;
      default: n3298_o = n2171_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1921:49  */
  always @*
    case (n3282_o)
      5'b10000: n3299_o = n3184_o;
      5'b01000: n3299_o = n3184_o;
      5'b00100: n3299_o = n3184_o;
      5'b00010: n3299_o = n3184_o;
      5'b00001: n3299_o = 1'b1;
      default: n3299_o = n3184_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1921:49  */
  always @*
    case (n3282_o)
      5'b10000: n3303_o = n3279_o;
      5'b01000: n3303_o = 7'b0010011;
      5'b00100: n3303_o = 7'b0000111;
      5'b00010: n3303_o = 7'b0000001;
      5'b00001: n3303_o = n2180_o;
      default: n3303_o = n2180_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3304_o = n3315_o ? n3284_o : n2026_o;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3305_o = n3316_o ? n3286_o : n2151_o;
  assign n3306_o = {n3296_o, n3292_o};
  assign n3307_o = n1909_o[40];
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3308_o = n3337_o ? n3288_o : n3307_o;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3309_o = n3338_o ? n3306_o : n2166_o;
  /* TG68KdotC_Kernel.vhd:1920:41  */
  assign n3310_o = n3221_o ? n3297_o : n2168_o;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3311_o = n3342_o ? n3298_o : n2171_o;
  /* TG68KdotC_Kernel.vhd:1920:41  */
  assign n3312_o = n3221_o ? n3299_o : n3184_o;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3313_o = n3347_o ? n3303_o : n2180_o;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3314_o = n3166_o ? n3194_o : n1921_o;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3315_o = n3221_o & n3166_o;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3316_o = n3221_o & n3166_o;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3318_o = n3166_o ? n3198_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3321_o = n3166_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3323_o = n3166_o ? n3210_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3325_o = n3166_o ? n3213_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3328_o = n3166_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3331_o = n3166_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3334_o = n3166_o ? 1'b1 : 1'b0;
  assign n3335_o = {n3310_o, n3173_o};
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3337_o = n3221_o & n3166_o;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3338_o = n3221_o & n3166_o;
  assign n3339_o = n1909_o[49];
  assign n3340_o = {n2168_o, n3339_o};
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3341_o = n3166_o ? n3335_o : n3340_o;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3342_o = n3221_o & n3166_o;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3344_o = n3166_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3346_o = n3166_o ? n3312_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1890:33  */
  assign n3347_o = n3221_o & n3166_o;
  /* TG68KdotC_Kernel.vhd:1889:25  */
  assign n3349_o = n2185_o == 4'b0001;
  /* TG68KdotC_Kernel.vhd:1889:36  */
  assign n3351_o = n2185_o == 4'b0010;
  /* TG68KdotC_Kernel.vhd:1889:36  */
  assign n3352_o = n3349_o | n3351_o;
  /* TG68KdotC_Kernel.vhd:1889:43  */
  assign n3354_o = n2185_o == 4'b0011;
  /* TG68KdotC_Kernel.vhd:1889:43  */
  assign n3355_o = n3352_o | n3354_o;
  /* TG68KdotC_Kernel.vhd:1966:42  */
  assign n3356_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:1967:50  */
  assign n3357_o = opcode[6];
  /* TG68KdotC_Kernel.vhd:1968:58  */
  assign n3358_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:1968:71  */
  assign n3360_o = n3358_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:1968:88  */
  assign n3361_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1968:100  */
  assign n3363_o = n3361_o == 3'b000;
  /* TG68KdotC_Kernel.vhd:1968:78  */
  assign n3364_o = n3363_o & n3360_o;
  /* TG68KdotC_Kernel.vhd:1969:66  */
  assign n3365_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:1969:81  */
  assign n3366_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:1969:74  */
  assign n3367_o = n3366_o & n3365_o;
  /* TG68KdotC_Kernel.vhd:1969:57  */
  assign n3374_o = n3367_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1969:57  */
  assign n3377_o = n3367_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1969:57  */
  assign n3380_o = n3367_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1969:57  */
  assign n3382_o = n3367_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1969:57  */
  assign n3384_o = n3367_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1969:57  */
  assign n3386_o = n3367_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1969:57  */
  assign n3388_o = n3367_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1980:66  */
  assign n3389_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:1981:67  */
  assign n3390_o = opcode[5];
  /* TG68KdotC_Kernel.vhd:1981:84  */
  assign n3391_o = opcode[4:3];
  /* TG68KdotC_Kernel.vhd:1981:96  */
  assign n3393_o = n3391_o == 2'b10;
  /* TG68KdotC_Kernel.vhd:1981:75  */
  assign n3394_o = n3390_o | n3393_o;
  /* TG68KdotC_Kernel.vhd:1980:74  */
  assign n3395_o = n3394_o & n3389_o;
  /* TG68KdotC_Kernel.vhd:1982:66  */
  assign n3396_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1982:78  */
  assign n3398_o = n3396_o != 3'b100;
  /* TG68KdotC_Kernel.vhd:1981:103  */
  assign n3399_o = n3398_o & n3395_o;
  /* TG68KdotC_Kernel.vhd:1982:96  */
  assign n3400_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:1982:108  */
  assign n3402_o = n3400_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:1982:86  */
  assign n3403_o = n3402_o & n3399_o;
  /* TG68KdotC_Kernel.vhd:1989:74  */
  assign n3407_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:1989:86  */
  assign n3409_o = n3407_o == 3'b010;
  /* TG68KdotC_Kernel.vhd:1989:65  */
  assign n3412_o = n3409_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1989:65  */
  assign n3415_o = n3409_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1989:65  */
  assign n3418_o = n3409_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1995:71  */
  assign n3419_o = set[62];
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3421_o = n3428_o ? 2'b01 : n2026_o;
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3423_o = n3442_o ? 1'b1 : n2154_o;
  /* TG68KdotC_Kernel.vhd:1999:65  */
  assign n3425_o = setexecopc ? 1'b1 : n3412_o;
  /* TG68KdotC_Kernel.vhd:1999:65  */
  assign n3427_o = setexecopc ? 1'b1 : n3415_o;
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3428_o = n3419_o & n3403_o;
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3431_o = n3403_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3434_o = n3403_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3437_o = n3403_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3439_o = n3403_o ? n3425_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3441_o = n3403_o ? n3427_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3442_o = n3419_o & n3403_o;
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3445_o = n3403_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3448_o = n3403_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3450_o = n3403_o ? n3418_o : 1'b0;
  assign n3451_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3452_o = n3403_o ? 1'b1 : n3451_o;
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3454_o = n3403_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1980:57  */
  assign n3456_o = n3403_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3457_o = n3364_o ? n2026_o : n3421_o;
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3459_o = n3364_o ? 1'b0 : n3431_o;
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3461_o = n3364_o ? 1'b0 : n3434_o;
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3462_o = n3364_o ? n3374_o : n3437_o;
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3464_o = n3364_o ? 1'b0 : n3439_o;
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3466_o = n3364_o ? 1'b0 : n3441_o;
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3467_o = n3364_o ? n2154_o : n3423_o;
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3468_o = n3364_o ? n3377_o : n3445_o;
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3469_o = n3364_o ? n3380_o : n3448_o;
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3471_o = n3364_o ? 1'b0 : n3450_o;
  assign n3472_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3473_o = n3364_o ? n3472_o : n3452_o;
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3474_o = n3364_o ? n3382_o : n3454_o;
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3476_o = n3364_o ? n3384_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3477_o = n3364_o ? n3386_o : n3456_o;
  /* TG68KdotC_Kernel.vhd:1968:49  */
  assign n3479_o = n3364_o ? n3388_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2009:58  */
  assign n3480_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2009:70  */
  assign n3482_o = n3480_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2010:59  */
  assign n3483_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2010:71  */
  assign n3485_o = n3483_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2010:89  */
  assign n3486_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:2010:101  */
  assign n3488_o = n3486_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2010:80  */
  assign n3489_o = n3485_o | n3488_o;
  /* TG68KdotC_Kernel.vhd:2009:78  */
  assign n3490_o = n3489_o & n3482_o;
  /* TG68KdotC_Kernel.vhd:2011:66  */
  assign n3491_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:2014:74  */
  assign n3493_o = c_out[1];
  /* TG68KdotC_Kernel.vhd:2014:77  */
  assign n3494_o = ~n3493_o;
  /* TG68KdotC_Kernel.vhd:2014:91  */
  assign n3495_o = op1out[15];
  /* TG68KdotC_Kernel.vhd:2014:82  */
  assign n3496_o = n3494_o | n3495_o;
  /* TG68KdotC_Kernel.vhd:2014:109  */
  assign n3497_o = op2out[15];
  /* TG68KdotC_Kernel.vhd:2014:100  */
  assign n3498_o = n3496_o | n3497_o;
  /* TG68KdotC_Kernel.vhd:2014:127  */
  assign n3499_o = exec[31];
  /* TG68KdotC_Kernel.vhd:2014:119  */
  assign n3500_o = n3499_o & n3498_o;
  /* TG68KdotC_Kernel.vhd:2014:65  */
  assign n3503_o = n3500_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2017:66  */
  assign n3504_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:2020:74  */
  assign n3506_o = c_out[2];
  /* TG68KdotC_Kernel.vhd:2020:77  */
  assign n3507_o = ~n3506_o;
  /* TG68KdotC_Kernel.vhd:2020:91  */
  assign n3508_o = op1out[31];
  /* TG68KdotC_Kernel.vhd:2020:82  */
  assign n3509_o = n3507_o | n3508_o;
  /* TG68KdotC_Kernel.vhd:2020:109  */
  assign n3510_o = op2out[31];
  /* TG68KdotC_Kernel.vhd:2020:100  */
  assign n3511_o = n3509_o | n3510_o;
  /* TG68KdotC_Kernel.vhd:2020:127  */
  assign n3512_o = exec[31];
  /* TG68KdotC_Kernel.vhd:2020:119  */
  assign n3513_o = n3512_o & n3511_o;
  /* TG68KdotC_Kernel.vhd:2020:65  */
  assign n3516_o = n3513_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2017:57  */
  assign n3518_o = n3504_o ? 2'b10 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2017:57  */
  assign n3521_o = n3504_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2017:57  */
  assign n3523_o = n3504_o ? n3516_o : 1'b1;
  assign n3524_o = n1909_o[43];
  /* TG68KdotC_Kernel.vhd:2017:57  */
  assign n3525_o = n3504_o ? 1'b1 : n3524_o;
  /* TG68KdotC_Kernel.vhd:2011:57  */
  assign n3527_o = n3491_o ? 2'b01 : n3518_o;
  /* TG68KdotC_Kernel.vhd:2011:57  */
  assign n3529_o = n3491_o ? 1'b0 : n3521_o;
  /* TG68KdotC_Kernel.vhd:2011:57  */
  assign n3530_o = n3491_o ? n3503_o : n3523_o;
  /* TG68KdotC_Kernel.vhd:2011:57  */
  assign n3531_o = n3491_o ? 1'b1 : n3525_o;
  /* TG68KdotC_Kernel.vhd:2027:66  */
  assign n3532_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:2027:80  */
  assign n3533_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:2027:74  */
  assign n3534_o = n3532_o | n3533_o;
  /* TG68KdotC_Kernel.vhd:2028:91  */
  assign n3535_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2028:103  */
  assign n3537_o = n3535_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2028:82  */
  assign n3538_o = nextpass | n3537_o;
  /* TG68KdotC_Kernel.vhd:2028:118  */
  assign n3539_o = exec[31];
  /* TG68KdotC_Kernel.vhd:2028:126  */
  assign n3540_o = ~n3539_o;
  /* TG68KdotC_Kernel.vhd:2028:110  */
  assign n3541_o = n3540_o & n3538_o;
  /* TG68KdotC_Kernel.vhd:2028:146  */
  assign n3543_o = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:2028:131  */
  assign n3544_o = n3543_o & n3541_o;
  /* TG68KdotC_Kernel.vhd:2028:65  */
  assign n3547_o = n3544_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2033:65  */
  assign n3551_o = setexecopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2033:65  */
  assign n3554_o = setexecopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2027:57  */
  assign n3556_o = n3534_o ? n3551_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2027:57  */
  assign n3558_o = n3534_o ? n3554_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2027:57  */
  assign n3561_o = n3534_o ? 1'b1 : 1'b0;
  assign n3562_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2009:49  */
  assign n3563_o = n3580_o ? 1'b1 : n3562_o;
  /* TG68KdotC_Kernel.vhd:2027:57  */
  assign n3565_o = n3534_o ? n3547_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2009:49  */
  assign n3566_o = n3490_o ? n3527_o : n1921_o;
  /* TG68KdotC_Kernel.vhd:2009:49  */
  assign n3568_o = n3490_o ? n3556_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2009:49  */
  assign n3570_o = n3490_o ? n3558_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2009:49  */
  assign n3572_o = n3490_o ? n3529_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:2009:49  */
  assign n3574_o = n3490_o ? n3530_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:2009:49  */
  assign n3576_o = n3490_o ? n3561_o : 1'b0;
  assign n3577_o = n1909_o[43];
  /* TG68KdotC_Kernel.vhd:2009:49  */
  assign n3578_o = n3490_o ? n3531_o : n3577_o;
  /* TG68KdotC_Kernel.vhd:2009:49  */
  assign n3580_o = n3534_o & n3490_o;
  /* TG68KdotC_Kernel.vhd:2009:49  */
  assign n3582_o = n3490_o ? n3565_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3583_o = n3357_o ? n1921_o : n3566_o;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3584_o = n3357_o ? n3457_o : n2026_o;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3586_o = n3357_o ? n3459_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3588_o = n3357_o ? n3461_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3589_o = n3357_o ? n3462_o : n3568_o;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3591_o = n3357_o ? n3464_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3592_o = n3357_o ? n3466_o : n3570_o;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3593_o = n3357_o ? n3467_o : n2154_o;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3594_o = n3357_o ? n3468_o : n3572_o;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3595_o = n3357_o ? n3469_o : n3574_o;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3596_o = n3357_o ? n3471_o : n3576_o;
  assign n3597_o = n1909_o[43];
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3598_o = n3357_o ? n3597_o : n3578_o;
  assign n3599_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3600_o = n3357_o ? n3473_o : n3599_o;
  assign n3601_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3602_o = n3357_o ? n3601_o : n3563_o;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3604_o = n3357_o ? n3474_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3606_o = n3357_o ? n3476_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3608_o = n3357_o ? 1'b0 : n3582_o;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3610_o = n3357_o ? n3477_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1967:41  */
  assign n3612_o = n3357_o ? n3479_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2044:52  */
  assign n3613_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:2046:67  */
  assign n3614_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2046:79  */
  assign n3616_o = n3614_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2047:67  */
  assign n3617_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2047:79  */
  assign n3619_o = n3617_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:2047:96  */
  assign n3620_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2047:108  */
  assign n3622_o = n3620_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2047:87  */
  assign n3623_o = n3619_o | n3622_o;
  /* TG68KdotC_Kernel.vhd:2046:87  */
  assign n3624_o = n3623_o & n3616_o;
  /* TG68KdotC_Kernel.vhd:2048:74  */
  assign n3625_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2048:86  */
  assign n3627_o = n3625_o == 2'b11;
  /* TG68KdotC_Kernel.vhd:2054:87  */
  assign n3629_o = cpu[0];
  /* TG68KdotC_Kernel.vhd:2054:104  */
  assign n3631_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:2054:95  */
  assign n3632_o = n3631_o & n3629_o;
  /* TG68KdotC_Kernel.vhd:2054:123  */
  assign n3633_o = ~addrvalue;
  /* TG68KdotC_Kernel.vhd:2054:110  */
  assign n3634_o = n3633_o & n3632_o;
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3636_o = n3672_o ? 1'b1 : make_berr;
  /* TG68KdotC_Kernel.vhd:2057:90  */
  assign n3637_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2057:102  */
  assign n3639_o = n3637_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2057:81  */
  assign n3642_o = n3639_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2071:82  */
  assign n3646_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2071:94  */
  assign n3648_o = n3646_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2071:73  */
  assign n3651_o = n3648_o ? 1'b1 : 1'b0;
  assign n3653_o = n1909_o[54];
  /* TG68KdotC_Kernel.vhd:2074:73  */
  assign n3654_o = setexecopc ? 1'b1 : n3653_o;
  /* TG68KdotC_Kernel.vhd:2048:65  */
  assign n3655_o = n3634_o & n3627_o;
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3657_o = n3673_o ? 2'b01 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2048:65  */
  assign n3660_o = n3627_o ? 1'b0 : 1'b1;
  assign n3661_o = n1909_o[54];
  /* TG68KdotC_Kernel.vhd:2048:65  */
  assign n3662_o = n3627_o ? n3661_o : n3654_o;
  assign n3663_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2048:65  */
  assign n3664_o = n3627_o ? n3663_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:2048:65  */
  assign n3666_o = n3627_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2048:65  */
  assign n3668_o = n3627_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2048:65  */
  assign n3670_o = n3627_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2048:65  */
  assign n3671_o = n3627_o ? n3642_o : n3651_o;
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3672_o = n3655_o & n3624_o;
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3673_o = n3627_o & n3624_o;
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3676_o = n3624_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3678_o = n3624_o ? n3660_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3681_o = n3624_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3684_o = n3624_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3687_o = n3624_o ? 1'b1 : 1'b0;
  assign n3688_o = n1909_o[54];
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3689_o = n3624_o ? n3662_o : n3688_o;
  assign n3690_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3691_o = n3624_o ? n3664_o : n3690_o;
  assign n3692_o = {n3668_o, n3666_o};
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3694_o = n3624_o ? n3692_o : 2'b00;
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3696_o = n3624_o ? n3670_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2046:57  */
  assign n3698_o = n3624_o ? n3671_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2045:49  */
  assign n3700_o = n3613_o == 3'b000;
  /* TG68KdotC_Kernel.vhd:2083:67  */
  assign n3701_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2083:79  */
  assign n3703_o = n3701_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2084:67  */
  assign n3704_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2084:79  */
  assign n3706_o = n3704_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:2084:96  */
  assign n3707_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2084:108  */
  assign n3709_o = n3707_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2084:87  */
  assign n3710_o = n3706_o | n3709_o;
  /* TG68KdotC_Kernel.vhd:2083:87  */
  assign n3711_o = n3710_o & n3703_o;
  /* TG68KdotC_Kernel.vhd:2085:74  */
  assign n3712_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2085:86  */
  assign n3714_o = n3712_o == 2'b11;
  /* TG68KdotC_Kernel.vhd:2105:71  */
  assign n3717_o = cpu[0];
  /* TG68KdotC_Kernel.vhd:2105:88  */
  assign n3719_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:2105:79  */
  assign n3720_o = n3719_o & n3717_o;
  /* TG68KdotC_Kernel.vhd:2105:107  */
  assign n3721_o = ~addrvalue;
  /* TG68KdotC_Kernel.vhd:2105:94  */
  assign n3722_o = n3721_o & n3720_o;
  /* TG68KdotC_Kernel.vhd:2105:65  */
  assign n3724_o = n3722_o ? 1'b1 : make_berr;
  assign n3726_o = n1909_o[54];
  /* TG68KdotC_Kernel.vhd:2108:73  */
  assign n3727_o = setexecopc ? 1'b1 : n3726_o;
  /* TG68KdotC_Kernel.vhd:2111:82  */
  assign n3728_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2111:94  */
  assign n3730_o = n3728_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2111:73  */
  assign n3733_o = n3730_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2085:65  */
  assign n3734_o = n3714_o ? make_berr : n3724_o;
  /* TG68KdotC_Kernel.vhd:2085:65  */
  assign n3737_o = n3714_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2085:65  */
  assign n3740_o = n3714_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2085:65  */
  assign n3743_o = n3714_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2085:65  */
  assign n3746_o = n3714_o ? 1'b0 : 1'b1;
  assign n3747_o = n1909_o[54];
  /* TG68KdotC_Kernel.vhd:2085:65  */
  assign n3748_o = n3714_o ? n3747_o : n3727_o;
  /* TG68KdotC_Kernel.vhd:2085:65  */
  assign n3750_o = n3714_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2085:65  */
  assign n3752_o = n3714_o ? 1'b0 : n3733_o;
  /* TG68KdotC_Kernel.vhd:2083:57  */
  assign n3753_o = n3711_o ? n3734_o : make_berr;
  /* TG68KdotC_Kernel.vhd:2083:57  */
  assign n3755_o = n3711_o ? n3737_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2083:57  */
  assign n3757_o = n3711_o ? n3740_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:2083:57  */
  assign n3759_o = n3711_o ? n3743_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:2083:57  */
  assign n3761_o = n3711_o ? n3746_o : 1'b0;
  assign n3762_o = n1909_o[54];
  /* TG68KdotC_Kernel.vhd:2083:57  */
  assign n3763_o = n3711_o ? n3748_o : n3762_o;
  /* TG68KdotC_Kernel.vhd:2083:57  */
  assign n3765_o = n3711_o ? n3750_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2083:57  */
  assign n3767_o = n3711_o ? n3752_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2082:49  */
  assign n3769_o = n3613_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:2120:66  */
  assign n3770_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2120:78  */
  assign n3772_o = n3770_o == 2'b11;
  /* TG68KdotC_Kernel.vhd:2121:74  */
  assign n3773_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2121:86  */
  assign n3775_o = n3773_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2122:75  */
  assign n3776_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2122:87  */
  assign n3778_o = n3776_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2122:105  */
  assign n3779_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:2122:117  */
  assign n3781_o = n3779_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2122:96  */
  assign n3782_o = n3778_o | n3781_o;
  /* TG68KdotC_Kernel.vhd:2121:94  */
  assign n3783_o = n3782_o & n3775_o;
  /* TG68KdotC_Kernel.vhd:2126:101  */
  assign n3784_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2126:113  */
  assign n3786_o = n3784_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2126:91  */
  assign n3787_o = n3786_o & decodeopc;
  /* TG68KdotC_Kernel.vhd:2126:129  */
  assign n3789_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:2126:148  */
  assign n3790_o = ~addrvalue;
  /* TG68KdotC_Kernel.vhd:2126:135  */
  assign n3791_o = n3790_o & n3789_o;
  /* TG68KdotC_Kernel.vhd:2126:120  */
  assign n3792_o = n3787_o | n3791_o;
  /* TG68KdotC_Kernel.vhd:2126:154  */
  assign n3793_o = n3792_o | direct_data;
  assign n3795_o = n1909_o[51];
  /* TG68KdotC_Kernel.vhd:2120:57  */
  assign n3796_o = n3866_o ? 1'b1 : n3795_o;
  /* TG68KdotC_Kernel.vhd:2120:57  */
  assign n3798_o = n3858_o ? 2'b01 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2121:65  */
  assign n3801_o = n3783_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2121:65  */
  assign n3804_o = n3783_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2121:65  */
  assign n3807_o = n3783_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2121:65  */
  assign n3810_o = n3783_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2121:65  */
  assign n3812_o = n3793_o & n3783_o;
  /* TG68KdotC_Kernel.vhd:2134:75  */
  assign n3813_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2134:87  */
  assign n3815_o = n3813_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2135:75  */
  assign n3816_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2135:87  */
  assign n3818_o = n3816_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:2135:104  */
  assign n3819_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2135:116  */
  assign n3821_o = n3819_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2135:95  */
  assign n3822_o = n3818_o | n3821_o;
  /* TG68KdotC_Kernel.vhd:2134:95  */
  assign n3823_o = n3822_o & n3815_o;
  /* TG68KdotC_Kernel.vhd:2141:82  */
  assign n3826_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2141:94  */
  assign n3828_o = n3826_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2141:73  */
  assign n3831_o = n3828_o ? 1'b1 : 1'b0;
  assign n3833_o = n1909_o[54];
  /* TG68KdotC_Kernel.vhd:2134:65  */
  assign n3834_o = n3851_o ? 1'b1 : n3833_o;
  /* TG68KdotC_Kernel.vhd:2134:65  */
  assign n3837_o = n3823_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2134:65  */
  assign n3840_o = n3823_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2134:65  */
  assign n3843_o = n3823_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2134:65  */
  assign n3846_o = n3823_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2134:65  */
  assign n3849_o = n3823_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2134:65  */
  assign n3851_o = setexecopc & n3823_o;
  assign n3852_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2134:65  */
  assign n3853_o = n3823_o ? 1'b1 : n3852_o;
  /* TG68KdotC_Kernel.vhd:2134:65  */
  assign n3855_o = n3823_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2134:65  */
  assign n3857_o = n3823_o ? n3831_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2120:57  */
  assign n3858_o = n3783_o & n3772_o;
  /* TG68KdotC_Kernel.vhd:2120:57  */
  assign n3860_o = n3772_o ? 1'b0 : n3837_o;
  /* TG68KdotC_Kernel.vhd:2120:57  */
  assign n3861_o = n3772_o ? n3801_o : n3840_o;
  /* TG68KdotC_Kernel.vhd:2120:57  */
  assign n3862_o = n3772_o ? n3804_o : n3843_o;
  /* TG68KdotC_Kernel.vhd:2120:57  */
  assign n3863_o = n3772_o ? n3807_o : n3846_o;
  /* TG68KdotC_Kernel.vhd:2120:57  */
  assign n3864_o = n3772_o ? n3810_o : n3849_o;
  /* TG68KdotC_Kernel.vhd:2120:57  */
  assign n3866_o = n3812_o & n3772_o;
  assign n3867_o = n1909_o[54];
  /* TG68KdotC_Kernel.vhd:2120:57  */
  assign n3868_o = n3772_o ? n3867_o : n3834_o;
  assign n3869_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2120:57  */
  assign n3870_o = n3772_o ? n3869_o : n3853_o;
  /* TG68KdotC_Kernel.vhd:2120:57  */
  assign n3872_o = n3772_o ? 1'b0 : n3855_o;
  /* TG68KdotC_Kernel.vhd:2120:57  */
  assign n3874_o = n3772_o ? 1'b0 : n3857_o;
  /* TG68KdotC_Kernel.vhd:2119:49  */
  assign n3876_o = n3613_o == 3'b010;
  /* TG68KdotC_Kernel.vhd:2153:66  */
  assign n3877_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2153:78  */
  assign n3879_o = n3877_o == 2'b11;
  /* TG68KdotC_Kernel.vhd:2154:74  */
  assign n3880_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2154:86  */
  assign n3882_o = n3880_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2155:75  */
  assign n3883_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2155:87  */
  assign n3885_o = n3883_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2155:105  */
  assign n3886_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:2155:117  */
  assign n3888_o = n3886_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2155:96  */
  assign n3889_o = n3885_o | n3888_o;
  /* TG68KdotC_Kernel.vhd:2154:94  */
  assign n3890_o = n3889_o & n3882_o;
  /* TG68KdotC_Kernel.vhd:2160:109  */
  assign n3891_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2160:121  */
  assign n3893_o = n3891_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2160:99  */
  assign n3894_o = n3893_o & decodeopc;
  /* TG68KdotC_Kernel.vhd:2160:137  */
  assign n3896_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:2160:156  */
  assign n3897_o = ~addrvalue;
  /* TG68KdotC_Kernel.vhd:2160:143  */
  assign n3898_o = n3897_o & n3896_o;
  /* TG68KdotC_Kernel.vhd:2160:128  */
  assign n3899_o = n3894_o | n3898_o;
  /* TG68KdotC_Kernel.vhd:2160:162  */
  assign n3900_o = n3899_o | direct_data;
  assign n3903_o = {1'b1, 1'b1};
  assign n3904_o = n1909_o[52:51];
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n3905_o = n4006_o ? n3903_o : n3904_o;
  /* TG68KdotC_Kernel.vhd:2164:88  */
  assign n3906_o = exec[52];
  /* TG68KdotC_Kernel.vhd:2164:128  */
  assign n3907_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2164:140  */
  assign n3909_o = n3907_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2164:118  */
  assign n3910_o = n3909_o & decodeopc;
  /* TG68KdotC_Kernel.vhd:2164:100  */
  assign n3911_o = n3906_o | n3910_o;
  /* TG68KdotC_Kernel.vhd:2164:156  */
  assign n3913_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:2164:175  */
  assign n3914_o = ~addrvalue;
  /* TG68KdotC_Kernel.vhd:2164:162  */
  assign n3915_o = n3914_o & n3913_o;
  /* TG68KdotC_Kernel.vhd:2164:147  */
  assign n3916_o = n3911_o | n3915_o;
  /* TG68KdotC_Kernel.vhd:2164:181  */
  assign n3917_o = n3916_o | direct_data;
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n3919_o = n3995_o ? 2'b01 : n2026_o;
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n3921_o = n3994_o ? 2'b01 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2156:73  */
  assign n3922_o = n3917_o & svmode;
  /* TG68KdotC_Kernel.vhd:2156:73  */
  assign n3925_o = svmode ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2156:73  */
  assign n3928_o = svmode ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2156:73  */
  assign n3931_o = svmode ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2156:73  */
  assign n3934_o = svmode ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2156:73  */
  assign n3936_o = n3900_o & svmode;
  /* TG68KdotC_Kernel.vhd:2154:65  */
  assign n3937_o = svmode & n3890_o;
  /* TG68KdotC_Kernel.vhd:2154:65  */
  assign n3938_o = n3922_o & n3890_o;
  /* TG68KdotC_Kernel.vhd:2154:65  */
  assign n3940_o = n3890_o ? n3925_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2154:65  */
  assign n3943_o = n3890_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2154:65  */
  assign n3945_o = n3890_o ? n3928_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2154:65  */
  assign n3947_o = n3890_o ? n3931_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:2154:65  */
  assign n3949_o = n3890_o ? n3934_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2154:65  */
  assign n3951_o = n3936_o & n3890_o;
  /* TG68KdotC_Kernel.vhd:2176:74  */
  assign n3952_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2176:86  */
  assign n3954_o = n3952_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2177:75  */
  assign n3955_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2177:87  */
  assign n3957_o = n3955_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:2177:104  */
  assign n3958_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2177:116  */
  assign n3960_o = n3958_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2177:95  */
  assign n3961_o = n3957_o | n3960_o;
  /* TG68KdotC_Kernel.vhd:2176:94  */
  assign n3962_o = n3961_o & n3954_o;
  /* TG68KdotC_Kernel.vhd:2182:82  */
  assign n3965_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2182:94  */
  assign n3967_o = n3965_o == 3'b000;
  /* TG68KdotC_Kernel.vhd:2182:73  */
  assign n3970_o = n3967_o ? 1'b1 : 1'b0;
  assign n3972_o = n1909_o[53];
  /* TG68KdotC_Kernel.vhd:2176:65  */
  assign n3973_o = n3987_o ? 1'b1 : n3972_o;
  /* TG68KdotC_Kernel.vhd:2176:65  */
  assign n3976_o = n3962_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2176:65  */
  assign n3979_o = n3962_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2176:65  */
  assign n3982_o = n3962_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2176:65  */
  assign n3985_o = n3962_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2176:65  */
  assign n3987_o = setexecopc & n3962_o;
  /* TG68KdotC_Kernel.vhd:2176:65  */
  assign n3989_o = n3962_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2176:65  */
  assign n3991_o = n3962_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2176:65  */
  assign n3993_o = n3962_o ? n3970_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n3994_o = n3937_o & n3879_o;
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n3995_o = n3938_o & n3879_o;
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n3997_o = n3879_o ? 1'b0 : n3976_o;
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n3999_o = n3879_o ? n3940_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n4000_o = n3879_o ? n3943_o : n3979_o;
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n4002_o = n3879_o ? n3945_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n4003_o = n3879_o ? n3947_o : n3982_o;
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n4004_o = n3879_o ? n3949_o : n3985_o;
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n4006_o = n3951_o & n3879_o;
  assign n4007_o = n1909_o[53];
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n4008_o = n3879_o ? n4007_o : n3973_o;
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n4010_o = n3879_o ? 1'b0 : n3989_o;
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n4012_o = n3879_o ? 1'b0 : n3991_o;
  /* TG68KdotC_Kernel.vhd:2153:57  */
  assign n4014_o = n3879_o ? 1'b0 : n3993_o;
  /* TG68KdotC_Kernel.vhd:2152:49  */
  assign n4016_o = n3613_o == 3'b011;
  /* TG68KdotC_Kernel.vhd:2194:66  */
  assign n4017_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:2195:74  */
  assign n4018_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2195:86  */
  assign n4020_o = n4018_o == 3'b000;
  /* TG68KdotC_Kernel.vhd:2195:103  */
  assign n4021_o = opcode[10];
  /* TG68KdotC_Kernel.vhd:2195:107  */
  assign n4022_o = ~n4021_o;
  /* TG68KdotC_Kernel.vhd:2195:93  */
  assign n4023_o = n4022_o & n4020_o;
  /* TG68KdotC_Kernel.vhd:2200:82  */
  assign n4027_o = opcode[6];
  /* TG68KdotC_Kernel.vhd:2200:85  */
  assign n4028_o = ~n4027_o;
  /* TG68KdotC_Kernel.vhd:2200:73  */
  assign n4031_o = n4028_o ? 2'b01 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2200:73  */
  assign n4033_o = n4028_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2206:83  */
  assign n4034_o = opcode[10];
  /* TG68KdotC_Kernel.vhd:2206:103  */
  assign n4035_o = opcode[5];
  /* TG68KdotC_Kernel.vhd:2206:120  */
  assign n4036_o = opcode[4:3];
  /* TG68KdotC_Kernel.vhd:2206:132  */
  assign n4038_o = n4036_o == 2'b10;
  /* TG68KdotC_Kernel.vhd:2206:111  */
  assign n4039_o = n4035_o | n4038_o;
  /* TG68KdotC_Kernel.vhd:2207:83  */
  assign n4040_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2207:95  */
  assign n4042_o = n4040_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:2207:112  */
  assign n4043_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2207:124  */
  assign n4045_o = n4043_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2207:103  */
  assign n4046_o = n4042_o | n4045_o;
  /* TG68KdotC_Kernel.vhd:2206:139  */
  assign n4047_o = n4046_o & n4039_o;
  /* TG68KdotC_Kernel.vhd:2206:92  */
  assign n4048_o = n4034_o | n4047_o;
  /* TG68KdotC_Kernel.vhd:2208:83  */
  assign n4049_o = opcode[10];
  /* TG68KdotC_Kernel.vhd:2208:87  */
  assign n4050_o = ~n4049_o;
  /* TG68KdotC_Kernel.vhd:2208:102  */
  assign n4051_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2208:114  */
  assign n4053_o = n4051_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:2209:82  */
  assign n4054_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2209:94  */
  assign n4056_o = n4054_o != 3'b100;
  /* TG68KdotC_Kernel.vhd:2208:121  */
  assign n4057_o = n4056_o & n4053_o;
  /* TG68KdotC_Kernel.vhd:2210:82  */
  assign n4058_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2210:94  */
  assign n4060_o = n4058_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2209:102  */
  assign n4061_o = n4060_o & n4057_o;
  /* TG68KdotC_Kernel.vhd:2208:92  */
  assign n4062_o = n4050_o | n4061_o;
  /* TG68KdotC_Kernel.vhd:2207:133  */
  assign n4063_o = n4062_o & n4048_o;
  /* TG68KdotC_Kernel.vhd:2213:90  */
  assign n4065_o = opcode[6];
  /* TG68KdotC_Kernel.vhd:2213:93  */
  assign n4066_o = ~n4065_o;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4068_o = n4156_o ? 2'b01 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2216:91  */
  assign n4069_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2216:103  */
  assign n4071_o = n4069_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:2216:119  */
  assign n4072_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2216:131  */
  assign n4074_o = n4072_o == 3'b011;
  /* TG68KdotC_Kernel.vhd:2216:110  */
  assign n4075_o = n4071_o | n4074_o;
  /* TG68KdotC_Kernel.vhd:2216:148  */
  assign n4077_o = state == 2'b01;
  /* TG68KdotC_Kernel.vhd:2216:139  */
  assign n4078_o = n4077_o & n4075_o;
  /* TG68KdotC_Kernel.vhd:2216:81  */
  assign n4082_o = n4078_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2216:81  */
  assign n4084_o = n4078_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2220:90  */
  assign n4085_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2220:102  */
  assign n4087_o = n4085_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:2220:81  */
  assign n4091_o = n4087_o ? 1'b1 : 1'b0;
  assign n4092_o = n1909_o[48];
  /* TG68KdotC_Kernel.vhd:2220:81  */
  assign n4093_o = n4087_o ? 1'b1 : n4092_o;
  /* TG68KdotC_Kernel.vhd:2224:89  */
  assign n4095_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:2224:108  */
  assign n4096_o = ~addrvalue;
  /* TG68KdotC_Kernel.vhd:2224:95  */
  assign n4097_o = n4096_o & n4095_o;
  assign n4100_o = n1909_o[0];
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4101_o = n4171_o ? 1'b1 : n4100_o;
  assign n4102_o = n1909_o[34];
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4103_o = n4173_o ? 1'b1 : n4102_o;
  /* TG68KdotC_Kernel.vhd:2230:98  */
  assign n4105_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2230:110  */
  assign n4107_o = n4105_o == 3'b010;
  /* TG68KdotC_Kernel.vhd:2230:126  */
  assign n4108_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2230:138  */
  assign n4110_o = n4108_o == 3'b011;
  /* TG68KdotC_Kernel.vhd:2230:117  */
  assign n4111_o = n4107_o | n4110_o;
  /* TG68KdotC_Kernel.vhd:2230:154  */
  assign n4112_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2230:166  */
  assign n4114_o = n4112_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:2230:145  */
  assign n4115_o = n4111_o | n4114_o;
  assign n4117_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:2230:89  */
  assign n4118_o = n4115_o ? n4117_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:2230:89  */
  assign n4121_o = n4115_o ? 7'b0011010 : 7'b0000001;
  assign n4122_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4123_o = n4177_o ? n4118_o : n4122_o;
  assign n4124_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4125_o = n4184_o ? 1'b1 : n4124_o;
  /* TG68KdotC_Kernel.vhd:2228:81  */
  assign n4126_o = decodeopc ? n4121_o : n2180_o;
  /* TG68KdotC_Kernel.vhd:2237:87  */
  assign n4127_o = set[62];
  /* TG68KdotC_Kernel.vhd:2240:106  */
  assign n4129_o = opcode[10];
  /* TG68KdotC_Kernel.vhd:2240:110  */
  assign n4130_o = ~n4129_o;
  /* TG68KdotC_Kernel.vhd:2240:97  */
  assign n4134_o = n4130_o ? 2'b11 : 2'b10;
  assign n4135_o = n1909_o[40];
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4136_o = n4175_o ? 1'b1 : n4135_o;
  /* TG68KdotC_Kernel.vhd:2238:89  */
  assign n4139_o = movem_run ? n4134_o : 2'b01;
  /* TG68KdotC_Kernel.vhd:2238:89  */
  assign n4141_o = n4130_o & movem_run;
  assign n4142_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4143_o = n4180_o ? 1'b1 : n4142_o;
  assign n4144_o = n1909_o[69];
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4145_o = n4182_o ? 1'b1 : n4144_o;
  /* TG68KdotC_Kernel.vhd:2237:81  */
  assign n4147_o = n4155_o ? 7'b0011011 : n4126_o;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4148_o = n4157_o ? n4139_o : n2026_o;
  /* TG68KdotC_Kernel.vhd:2237:81  */
  assign n4150_o = n4141_o & n4127_o;
  /* TG68KdotC_Kernel.vhd:2237:81  */
  assign n4152_o = movem_run & n4127_o;
  /* TG68KdotC_Kernel.vhd:2237:81  */
  assign n4154_o = movem_run & n4127_o;
  /* TG68KdotC_Kernel.vhd:2237:81  */
  assign n4155_o = movem_run & n4127_o;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4156_o = n4066_o & n4063_o;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4157_o = n4127_o & n4063_o;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4160_o = n4063_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4162_o = n4063_o ? n4091_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4165_o = n4063_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4168_o = n4063_o ? 1'b0 : 1'b1;
  assign n4169_o = {1'b1, n4093_o};
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4171_o = n4097_o & n4063_o;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4173_o = n4097_o & n4063_o;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4175_o = n4150_o & n4063_o;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4177_o = decodeopc & n4063_o;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4178_o = n4063_o ? n4169_o : n2177_o;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4180_o = n4152_o & n4063_o;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4182_o = n4154_o & n4063_o;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4184_o = decodeopc & n4063_o;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4186_o = n4063_o ? n4082_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4188_o = n4063_o ? n4084_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2206:73  */
  assign n4189_o = n4063_o ? n4147_o : n2180_o;
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4190_o = n4023_o ? n4031_o : n4068_o;
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4191_o = n4023_o ? n2026_o : n4148_o;
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4193_o = n4023_o ? 1'b0 : n4160_o;
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4196_o = n4023_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4198_o = n4023_o ? 1'b0 : n4162_o;
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4200_o = n4023_o ? 1'b0 : n4165_o;
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4202_o = n4023_o ? 1'b0 : n4168_o;
  assign n4203_o = n1909_o[0];
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4204_o = n4023_o ? n4203_o : n4101_o;
  assign n4205_o = n1909_o[34];
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4206_o = n4023_o ? n4205_o : n4103_o;
  assign n4207_o = n1909_o[40];
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4208_o = n4023_o ? n4207_o : n4136_o;
  assign n4209_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4210_o = n4023_o ? n4209_o : n4123_o;
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4211_o = n4023_o ? n2177_o : n4178_o;
  assign n4212_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4213_o = n4023_o ? n4212_o : n4143_o;
  assign n4214_o = n1909_o[69];
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4215_o = n4023_o ? n4214_o : n4145_o;
  assign n4216_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4217_o = n4023_o ? n4216_o : n4125_o;
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4219_o = n4023_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4221_o = n4023_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4223_o = n4023_o ? 1'b0 : n4186_o;
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4224_o = n4023_o ? 1'b1 : n4188_o;
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4226_o = n4023_o ? n4033_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2195:65  */
  assign n4227_o = n4023_o ? n2180_o : n4189_o;
  /* TG68KdotC_Kernel.vhd:2258:74  */
  assign n4228_o = opcode[10];
  /* TG68KdotC_Kernel.vhd:2282:85  */
  assign n4244_o = opcode[8:7];
  /* TG68KdotC_Kernel.vhd:2282:97  */
  assign n4246_o = n4244_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2282:113  */
  assign n4247_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2282:125  */
  assign n4249_o = n4247_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2282:103  */
  assign n4250_o = n4249_o & n4246_o;
  /* TG68KdotC_Kernel.vhd:2282:144  */
  assign n4251_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2282:156  */
  assign n4253_o = n4251_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2282:174  */
  assign n4254_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:2282:186  */
  assign n4256_o = n4254_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2282:165  */
  assign n4257_o = n4253_o | n4256_o;
  /* TG68KdotC_Kernel.vhd:2282:133  */
  assign n4258_o = n4257_o & n4250_o;
  /* TG68KdotC_Kernel.vhd:2283:84  */
  assign n4259_o = opcode[6];
  /* TG68KdotC_Kernel.vhd:2283:115  */
  assign n4260_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:2283:123  */
  assign n4262_o = 1'b1 & n4260_o;
  /* TG68KdotC_Kernel.vhd:2283:108  */
  assign n4264_o = 1'b0 | n4262_o;
  /* TG68KdotC_Kernel.vhd:2283:92  */
  assign n4265_o = n4264_o & n4259_o;
  /* TG68KdotC_Kernel.vhd:2284:83  */
  assign n4266_o = opcode[6];
  /* TG68KdotC_Kernel.vhd:2284:86  */
  assign n4267_o = ~n4266_o;
  /* TG68KdotC_Kernel.vhd:2284:114  */
  assign n4268_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:2284:122  */
  assign n4270_o = 1'b1 & n4268_o;
  /* TG68KdotC_Kernel.vhd:2284:107  */
  assign n4272_o = 1'b0 | n4270_o;
  /* TG68KdotC_Kernel.vhd:2284:91  */
  assign n4273_o = n4272_o & n4267_o;
  /* TG68KdotC_Kernel.vhd:2283:141  */
  assign n4274_o = n4265_o | n4273_o;
  /* TG68KdotC_Kernel.vhd:2282:193  */
  assign n4275_o = n4274_o & n4258_o;
  assign n4278_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4279_o = n4618_o ? 1'b1 : n4278_o;
  assign n4280_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4281_o = n4630_o ? 1'b1 : n4280_o;
  /* TG68KdotC_Kernel.vhd:2285:81  */
  assign n4283_o = decodeopc ? 7'b0000001 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2290:96  */
  assign n4285_o = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:2290:102  */
  assign n4286_o = nextpass & n4285_o;
  /* TG68KdotC_Kernel.vhd:2290:130  */
  assign n4287_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2290:142  */
  assign n4289_o = n4287_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2290:156  */
  assign n4290_o = exec[42];
  /* TG68KdotC_Kernel.vhd:2290:148  */
  assign n4291_o = n4290_o & n4289_o;
  /* TG68KdotC_Kernel.vhd:2290:120  */
  assign n4292_o = n4286_o | n4291_o;
  /* TG68KdotC_Kernel.vhd:2294:98  */
  assign n4293_o = opcode[6];
  assign n4295_o = n1909_o[24];
  /* TG68KdotC_Kernel.vhd:2294:89  */
  assign n4296_o = n4293_o ? n4295_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:2294:89  */
  assign n4299_o = n4293_o ? 7'b1011001 : 7'b1010101;
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4301_o = n4321_o ? 2'b01 : n2026_o;
  /* TG68KdotC_Kernel.vhd:2290:81  */
  assign n4304_o = n4292_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2290:81  */
  assign n4307_o = n4292_o ? 1'b1 : 1'b0;
  assign n4308_o = n1909_o[24];
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4309_o = n4614_o ? n4296_o : n4308_o;
  /* TG68KdotC_Kernel.vhd:2290:81  */
  assign n4310_o = n4292_o ? n4299_o : n4283_o;
  /* TG68KdotC_Kernel.vhd:2302:107  */
  assign n4311_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2302:119  */
  assign n4313_o = n4311_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2302:125  */
  assign n4314_o = decodeopc & n4313_o;
  /* TG68KdotC_Kernel.vhd:2302:97  */
  assign n4315_o = nextpass | n4314_o;
  /* TG68KdotC_Kernel.vhd:2302:81  */
  assign n4318_o = n4315_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4320_o = n4275_o ? 2'b10 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4321_o = n4292_o & n4275_o;
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4324_o = n4275_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4326_o = n4275_o ? n4304_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4328_o = n4275_o ? n4307_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4330_o = n4275_o ? n4318_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4333_o = n4275_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4336_o = n4275_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4338_o = n4292_o & n4275_o;
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4340_o = decodeopc & n4275_o;
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4342_o = decodeopc & n4275_o;
  /* TG68KdotC_Kernel.vhd:2282:73  */
  assign n4343_o = n4275_o ? n4310_o : n2180_o;
  /* TG68KdotC_Kernel.vhd:2312:82  */
  assign n4344_o = opcode[6];
  /* TG68KdotC_Kernel.vhd:2314:90  */
  assign n4345_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2314:102  */
  assign n4347_o = n4345_o == 3'b000;
  /* TG68KdotC_Kernel.vhd:2317:93  */
  assign n4350_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2317:105  */
  assign n4352_o = n4350_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:2321:99  */
  assign n4353_o = opcode[5];
  /* TG68KdotC_Kernel.vhd:2321:116  */
  assign n4354_o = opcode[4:3];
  /* TG68KdotC_Kernel.vhd:2321:128  */
  assign n4356_o = n4354_o == 2'b10;
  /* TG68KdotC_Kernel.vhd:2321:107  */
  assign n4357_o = n4353_o | n4356_o;
  /* TG68KdotC_Kernel.vhd:2322:98  */
  assign n4358_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2322:110  */
  assign n4360_o = n4358_o != 3'b100;
  /* TG68KdotC_Kernel.vhd:2321:135  */
  assign n4361_o = n4360_o & n4357_o;
  /* TG68KdotC_Kernel.vhd:2323:98  */
  assign n4362_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2323:110  */
  assign n4364_o = n4362_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2322:118  */
  assign n4365_o = n4364_o & n4361_o;
  /* TG68KdotC_Kernel.vhd:2326:128  */
  assign n4367_o = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:2326:113  */
  assign n4368_o = n4367_o & nextpass;
  /* TG68KdotC_Kernel.vhd:2326:97  */
  assign n4371_o = n4368_o ? 2'b11 : n2026_o;
  /* TG68KdotC_Kernel.vhd:2321:89  */
  assign n4373_o = n4384_o ? 1'b1 : n2015_o;
  assign n4374_o = n2162_o[1];
  assign n4375_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n4376_o = n2037_o ? n4374_o : n4375_o;
  /* TG68KdotC_Kernel.vhd:2326:97  */
  assign n4377_o = n4368_o ? 1'b1 : n4376_o;
  /* TG68KdotC_Kernel.vhd:2321:89  */
  assign n4379_o = n4401_o ? 7'b0000001 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2332:103  */
  assign n4380_o = set[62];
  /* TG68KdotC_Kernel.vhd:2332:97  */
  assign n4382_o = n4380_o ? 2'b01 : n4371_o;
  /* TG68KdotC_Kernel.vhd:2321:89  */
  assign n4383_o = n4365_o ? n4382_o : n2026_o;
  /* TG68KdotC_Kernel.vhd:2321:89  */
  assign n4384_o = n4368_o & n4365_o;
  /* TG68KdotC_Kernel.vhd:2321:89  */
  assign n4387_o = n4365_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2321:89  */
  assign n4390_o = n4365_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2321:89  */
  assign n4393_o = n4365_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2321:89  */
  assign n4396_o = n4365_o ? 1'b1 : 1'b0;
  assign n4397_o = n2162_o[1];
  assign n4398_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n4399_o = n2037_o ? n4397_o : n4398_o;
  /* TG68KdotC_Kernel.vhd:2321:89  */
  assign n4400_o = n4365_o ? n4377_o : n4399_o;
  /* TG68KdotC_Kernel.vhd:2321:89  */
  assign n4401_o = n4368_o & n4365_o;
  /* TG68KdotC_Kernel.vhd:2317:81  */
  assign n4402_o = n4352_o ? n2026_o : n4383_o;
  /* TG68KdotC_Kernel.vhd:2317:81  */
  assign n4403_o = n4352_o ? n2015_o : n4373_o;
  /* TG68KdotC_Kernel.vhd:2317:81  */
  assign n4405_o = n4352_o ? 1'b0 : n4387_o;
  /* TG68KdotC_Kernel.vhd:2317:81  */
  assign n4407_o = n4352_o ? 1'b1 : n4390_o;
  /* TG68KdotC_Kernel.vhd:2317:81  */
  assign n4409_o = n4352_o ? 1'b1 : n4393_o;
  /* TG68KdotC_Kernel.vhd:2317:81  */
  assign n4411_o = n4352_o ? 1'b0 : n4396_o;
  assign n4412_o = n2162_o[1];
  assign n4413_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n4414_o = n2037_o ? n4412_o : n4413_o;
  /* TG68KdotC_Kernel.vhd:2317:81  */
  assign n4415_o = n4352_o ? n4414_o : n4400_o;
  /* TG68KdotC_Kernel.vhd:2317:81  */
  assign n4416_o = n4352_o ? n2180_o : n4379_o;
  /* TG68KdotC_Kernel.vhd:2314:81  */
  assign n4417_o = n4347_o ? n2026_o : n4402_o;
  /* TG68KdotC_Kernel.vhd:2314:81  */
  assign n4418_o = n4347_o ? n2015_o : n4403_o;
  /* TG68KdotC_Kernel.vhd:2314:81  */
  assign n4420_o = n4347_o ? 1'b0 : n4405_o;
  /* TG68KdotC_Kernel.vhd:2314:81  */
  assign n4422_o = n4347_o ? 1'b0 : n4407_o;
  /* TG68KdotC_Kernel.vhd:2314:81  */
  assign n4424_o = n4347_o ? 1'b0 : n4409_o;
  /* TG68KdotC_Kernel.vhd:2314:81  */
  assign n4426_o = n4347_o ? 1'b0 : n4411_o;
  assign n4427_o = n2162_o[1];
  assign n4428_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n4429_o = n2037_o ? n4427_o : n4428_o;
  /* TG68KdotC_Kernel.vhd:2314:81  */
  assign n4430_o = n4347_o ? n4429_o : n4415_o;
  /* TG68KdotC_Kernel.vhd:2314:81  */
  assign n4432_o = n4347_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2314:81  */
  assign n4434_o = n4347_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2314:81  */
  assign n4435_o = n4347_o ? n2180_o : n4416_o;
  /* TG68KdotC_Kernel.vhd:2341:90  */
  assign n4436_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2341:102  */
  assign n4438_o = n4436_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4448_o = n4523_o ? 1'b1 : n2015_o;
  /* TG68KdotC_Kernel.vhd:2346:89  */
  assign n4451_o = decodeopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2346:89  */
  assign n4454_o = decodeopc ? 1'b1 : 1'b0;
  assign n4455_o = n1909_o[36];
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4456_o = n4534_o ? 1'b1 : n4455_o;
  assign n4457_o = n1909_o[44];
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4458_o = n4536_o ? 1'b1 : n4457_o;
  assign n4459_o = n2162_o[1];
  assign n4460_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n4461_o = n2037_o ? n4459_o : n4460_o;
  /* TG68KdotC_Kernel.vhd:2346:89  */
  assign n4462_o = decodeopc ? 1'b1 : n4461_o;
  assign n4463_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4464_o = n4546_o ? 1'b1 : n4463_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4465_o = n4549_o ? 1'b1 : n2171_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4467_o = n4556_o ? 7'b0100011 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2358:98  */
  assign n4468_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2358:110  */
  assign n4470_o = n4468_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2359:99  */
  assign n4471_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2359:111  */
  assign n4473_o = n4471_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:2359:128  */
  assign n4474_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2359:140  */
  assign n4476_o = n4474_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2359:119  */
  assign n4477_o = n4473_o | n4476_o;
  /* TG68KdotC_Kernel.vhd:2358:118  */
  assign n4478_o = n4477_o & n4470_o;
  /* TG68KdotC_Kernel.vhd:2367:106  */
  assign n4483_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2367:118  */
  assign n4485_o = n4483_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2367:97  */
  assign n4488_o = n4485_o ? 1'b1 : 1'b0;
  assign n4490_o = n1909_o[54];
  /* TG68KdotC_Kernel.vhd:2358:89  */
  assign n4491_o = n4508_o ? 1'b1 : n4490_o;
  /* TG68KdotC_Kernel.vhd:2358:89  */
  assign n4494_o = n4478_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2358:89  */
  assign n4497_o = n4478_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2358:89  */
  assign n4500_o = n4478_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2358:89  */
  assign n4503_o = n4478_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2358:89  */
  assign n4506_o = n4478_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2358:89  */
  assign n4508_o = setexecopc & n4478_o;
  assign n4509_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2358:89  */
  assign n4510_o = n4478_o ? 1'b1 : n4509_o;
  /* TG68KdotC_Kernel.vhd:2358:89  */
  assign n4512_o = n4478_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2358:89  */
  assign n4514_o = n4478_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2358:89  */
  assign n4516_o = n4478_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2358:89  */
  assign n4518_o = n4478_o ? n4488_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4520_o = n4438_o ? 2'b10 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4522_o = n4438_o ? 1'b0 : n4494_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4523_o = decodeopc & n4438_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4525_o = n4438_o ? n4451_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4526_o = n4438_o ? n4454_o : n4497_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4528_o = n4438_o ? 1'b0 : n4500_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4530_o = n4438_o ? 1'b0 : n4503_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4532_o = n4438_o ? 1'b0 : n4506_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4534_o = decodeopc & n4438_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4536_o = decodeopc & n4438_o;
  assign n4537_o = n2162_o[1];
  assign n4538_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n4539_o = n2037_o ? n4537_o : n4538_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4540_o = n4438_o ? n4462_o : n4539_o;
  assign n4541_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4542_o = n4438_o ? 1'b1 : n4541_o;
  assign n4543_o = n1909_o[54];
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4544_o = n4438_o ? n4543_o : n4491_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4546_o = decodeopc & n4438_o;
  assign n4547_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4548_o = n4438_o ? n4547_o : n4510_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4549_o = decodeopc & n4438_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4550_o = n4438_o ? 1'b1 : n4512_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4552_o = n4438_o ? 1'b0 : n4514_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4554_o = n4438_o ? 1'b0 : n4516_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4555_o = n4438_o ? 1'b1 : n4518_o;
  /* TG68KdotC_Kernel.vhd:2341:81  */
  assign n4556_o = decodeopc & n4438_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4558_o = n4344_o ? 2'b10 : n4520_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4559_o = n4344_o ? n4417_o : n2026_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4561_o = n4344_o ? 1'b0 : n4522_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4562_o = n4344_o ? n4418_o : n4448_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4564_o = n4344_o ? n4420_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4566_o = n4344_o ? 1'b0 : n4525_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4568_o = n4344_o ? 1'b0 : n4526_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4569_o = n4344_o ? n4422_o : n4528_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4570_o = n4344_o ? n4424_o : n4530_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4571_o = n4344_o ? n4426_o : n4532_o;
  assign n4572_o = {n4548_o, n4464_o, n4544_o};
  assign n4573_o = n1909_o[36];
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4574_o = n4344_o ? n4573_o : n4456_o;
  assign n4575_o = n1909_o[44];
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4576_o = n4344_o ? n4575_o : n4458_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4577_o = n4344_o ? n4430_o : n4540_o;
  assign n4578_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4579_o = n4344_o ? n4578_o : n4542_o;
  assign n4580_o = n1909_o[56:54];
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4581_o = n4344_o ? n4580_o : n4572_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4582_o = n4344_o ? n2171_o : n4465_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4584_o = n4344_o ? 1'b0 : n4550_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4586_o = n4344_o ? 1'b0 : n4552_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4588_o = n4344_o ? n4432_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4590_o = n4344_o ? 1'b0 : n4554_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4591_o = n4344_o ? n4434_o : n4555_o;
  /* TG68KdotC_Kernel.vhd:2312:73  */
  assign n4592_o = n4344_o ? n4435_o : n4467_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4593_o = n4228_o ? n4320_o : n4558_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4594_o = n4228_o ? n4301_o : n4559_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4596_o = n4228_o ? 1'b0 : n4561_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4597_o = n4228_o ? n2015_o : n4562_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4599_o = n4228_o ? 1'b0 : n4564_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4601_o = n4228_o ? 1'b0 : n4566_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4602_o = n4228_o ? n4324_o : n4568_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4604_o = n4228_o ? n4326_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4606_o = n4228_o ? n4328_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4608_o = n4228_o ? n4330_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4609_o = n4228_o ? n4333_o : n4569_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4610_o = n4228_o ? n4336_o : n4570_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4612_o = n4228_o ? 1'b0 : n4571_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4614_o = n4338_o & n4228_o;
  assign n4615_o = n1909_o[36];
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4616_o = n4228_o ? n4615_o : n4574_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4618_o = n4340_o & n4228_o;
  assign n4619_o = n1909_o[44];
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4620_o = n4228_o ? n4619_o : n4576_o;
  assign n4621_o = n2162_o[1];
  assign n4622_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n4623_o = n2037_o ? n4621_o : n4622_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4624_o = n4228_o ? n4623_o : n4577_o;
  assign n4625_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4626_o = n4228_o ? n4625_o : n4579_o;
  assign n4627_o = n1909_o[56:54];
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4628_o = n4228_o ? n4627_o : n4581_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4630_o = n4342_o & n4228_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4631_o = n4228_o ? n2171_o : n4582_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4633_o = n4228_o ? 1'b0 : n4584_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4635_o = n4228_o ? 1'b0 : n4586_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4637_o = n4228_o ? 1'b0 : n4588_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4639_o = n4228_o ? 1'b0 : n4590_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4641_o = n4228_o ? 1'b0 : n4591_o;
  /* TG68KdotC_Kernel.vhd:2258:65  */
  assign n4642_o = n4228_o ? n4343_o : n4592_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4643_o = n4017_o ? n4190_o : n4593_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4644_o = n4017_o ? n4191_o : n4594_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4646_o = n4017_o ? 1'b0 : n4596_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4647_o = n4017_o ? n2015_o : n4597_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4648_o = n4017_o ? n4193_o : n4599_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4650_o = n4017_o ? 1'b0 : n4601_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4651_o = n4017_o ? n4196_o : n4602_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4653_o = n4017_o ? 1'b0 : n4604_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4655_o = n4017_o ? 1'b0 : n4606_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4657_o = n4017_o ? 1'b0 : n4608_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4659_o = n4017_o ? n4198_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4660_o = n4017_o ? n4200_o : n4609_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4661_o = n4017_o ? n4202_o : n4610_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4663_o = n4017_o ? 1'b0 : n4612_o;
  assign n4664_o = n1909_o[0];
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4665_o = n4017_o ? n4204_o : n4664_o;
  assign n4666_o = n1909_o[24];
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4667_o = n4017_o ? n4666_o : n4309_o;
  assign n4668_o = n1909_o[34];
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4669_o = n4017_o ? n4206_o : n4668_o;
  assign n4670_o = n1909_o[36];
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4671_o = n4017_o ? n4670_o : n4616_o;
  assign n4672_o = n1909_o[40];
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4673_o = n4017_o ? n4208_o : n4672_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4674_o = n4017_o ? n4210_o : n4279_o;
  assign n4675_o = n1909_o[44];
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4676_o = n4017_o ? n4675_o : n4620_o;
  assign n4677_o = n2162_o[1];
  assign n4678_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n4679_o = n2037_o ? n4677_o : n4678_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4680_o = n4017_o ? n4679_o : n4624_o;
  assign n4681_o = n4211_o[0];
  assign n4682_o = n1909_o[48];
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4683_o = n4017_o ? n4681_o : n4682_o;
  assign n4684_o = n4211_o[1];
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4685_o = n4017_o ? n4684_o : n4626_o;
  assign n4686_o = n4628_o[0];
  assign n4687_o = n1909_o[54];
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4688_o = n4017_o ? n4687_o : n4686_o;
  assign n4689_o = n4628_o[1];
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4690_o = n4017_o ? n4213_o : n4689_o;
  assign n4691_o = n4628_o[2];
  assign n4692_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4693_o = n4017_o ? n4692_o : n4691_o;
  assign n4694_o = n1909_o[69];
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4695_o = n4017_o ? n4215_o : n4694_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4696_o = n4017_o ? n4217_o : n4281_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4697_o = n4017_o ? n2171_o : n4631_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4699_o = n4017_o ? n4219_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4701_o = n4017_o ? 1'b0 : n4633_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4703_o = n4017_o ? n4221_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4705_o = n4017_o ? 1'b0 : n4635_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4707_o = n4017_o ? 1'b0 : n4637_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4709_o = n4017_o ? 1'b0 : n4639_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4711_o = n4017_o ? n4223_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4712_o = n4017_o ? n4224_o : n4641_o;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4714_o = n4017_o ? n4226_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2194:57  */
  assign n4715_o = n4017_o ? n4227_o : n4642_o;
  /* TG68KdotC_Kernel.vhd:2193:49  */
  assign n4717_o = n3613_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:2193:59  */
  assign n4719_o = n3613_o == 3'b110;
  /* TG68KdotC_Kernel.vhd:2193:59  */
  assign n4720_o = n4717_o | n4719_o;
  /* TG68KdotC_Kernel.vhd:2384:66  */
  assign n4721_o = opcode[7:3];
  /* TG68KdotC_Kernel.vhd:2384:78  */
  assign n4723_o = n4721_o == 5'b11111;
  /* TG68KdotC_Kernel.vhd:2384:97  */
  assign n4724_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2384:109  */
  assign n4726_o = n4724_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:2384:87  */
  assign n4727_o = n4726_o & n4723_o;
  /* TG68KdotC_Kernel.vhd:2388:75  */
  assign n4728_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2388:87  */
  assign n4730_o = n4728_o != 2'b11;
  /* TG68KdotC_Kernel.vhd:2389:75  */
  assign n4731_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2389:87  */
  assign n4733_o = n4731_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2390:75  */
  assign n4734_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2390:87  */
  assign n4736_o = n4734_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:2390:104  */
  assign n4737_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2390:116  */
  assign n4739_o = n4737_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2390:95  */
  assign n4740_o = n4736_o | n4739_o;
  /* TG68KdotC_Kernel.vhd:2389:95  */
  assign n4741_o = n4740_o & n4733_o;
  /* TG68KdotC_Kernel.vhd:2388:94  */
  assign n4742_o = n4730_o | n4741_o;
  /* TG68KdotC_Kernel.vhd:2391:76  */
  assign n4743_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2391:88  */
  assign n4745_o = n4743_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:2391:105  */
  assign n4746_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2391:117  */
  assign n4748_o = n4746_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2391:95  */
  assign n4749_o = n4745_o | n4748_o;
  /* TG68KdotC_Kernel.vhd:2392:75  */
  assign n4750_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2392:87  */
  assign n4752_o = n4750_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2392:105  */
  assign n4753_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:2392:117  */
  assign n4755_o = n4753_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2392:96  */
  assign n4756_o = n4752_o | n4755_o;
  /* TG68KdotC_Kernel.vhd:2391:127  */
  assign n4757_o = n4756_o & n4749_o;
  /* TG68KdotC_Kernel.vhd:2390:125  */
  assign n4758_o = n4757_o & n4742_o;
  /* TG68KdotC_Kernel.vhd:2396:90  */
  assign n4759_o = opcode[3];
  /* TG68KdotC_Kernel.vhd:2396:81  */
  assign n4762_o = n4759_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2394:73  */
  assign n4764_o = setexecopc ? n4762_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2394:73  */
  assign n4767_o = setexecopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2401:82  */
  assign n4769_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2401:94  */
  assign n4771_o = n4769_o == 2'b11;
  /* TG68KdotC_Kernel.vhd:2405:90  */
  assign n4772_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2405:102  */
  assign n4774_o = n4772_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2405:81  */
  assign n4777_o = n4774_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2388:65  */
  assign n4779_o = n4788_o ? 2'b00 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2401:73  */
  assign n4782_o = n4771_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2401:73  */
  assign n4785_o = n4771_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2401:73  */
  assign n4787_o = n4771_o ? n4777_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2388:65  */
  assign n4788_o = n4771_o & n4758_o;
  /* TG68KdotC_Kernel.vhd:2388:65  */
  assign n4790_o = n4758_o ? n4782_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2388:65  */
  assign n4792_o = n4758_o ? n4785_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2388:65  */
  assign n4794_o = n4758_o ? n4764_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2388:65  */
  assign n4796_o = n4758_o ? n4767_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2388:65  */
  assign n4799_o = n4758_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2388:65  */
  assign n4802_o = n4758_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2388:65  */
  assign n4805_o = n4758_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2388:65  */
  assign n4807_o = n4758_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2388:65  */
  assign n4809_o = n4758_o ? n4787_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2384:57  */
  assign n4810_o = n4727_o ? n1921_o : n4779_o;
  /* TG68KdotC_Kernel.vhd:2384:57  */
  assign n4812_o = n4727_o ? 1'b0 : n4790_o;
  /* TG68KdotC_Kernel.vhd:2384:57  */
  assign n4814_o = n4727_o ? 1'b0 : n4792_o;
  /* TG68KdotC_Kernel.vhd:2384:57  */
  assign n4816_o = n4727_o ? 1'b0 : n4794_o;
  /* TG68KdotC_Kernel.vhd:2384:57  */
  assign n4818_o = n4727_o ? 1'b0 : n4796_o;
  /* TG68KdotC_Kernel.vhd:2384:57  */
  assign n4820_o = n4727_o ? 1'b1 : n4799_o;
  /* TG68KdotC_Kernel.vhd:2384:57  */
  assign n4822_o = n4727_o ? 1'b1 : n4802_o;
  /* TG68KdotC_Kernel.vhd:2384:57  */
  assign n4824_o = n4727_o ? 1'b0 : n4805_o;
  /* TG68KdotC_Kernel.vhd:2384:57  */
  assign n4826_o = n4727_o ? 1'b0 : n4807_o;
  /* TG68KdotC_Kernel.vhd:2384:57  */
  assign n4828_o = n4727_o ? 1'b0 : n4809_o;
  /* TG68KdotC_Kernel.vhd:2382:49  */
  assign n4830_o = n3613_o == 3'b101;
  /* TG68KdotC_Kernel.vhd:2433:66  */
  assign n4831_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:2434:75  */
  assign n4832_o = opcode[5];
  /* TG68KdotC_Kernel.vhd:2434:92  */
  assign n4833_o = opcode[4:3];
  /* TG68KdotC_Kernel.vhd:2434:104  */
  assign n4835_o = n4833_o == 2'b10;
  /* TG68KdotC_Kernel.vhd:2434:83  */
  assign n4836_o = n4832_o | n4835_o;
  /* TG68KdotC_Kernel.vhd:2435:74  */
  assign n4837_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2435:86  */
  assign n4839_o = n4837_o != 3'b100;
  /* TG68KdotC_Kernel.vhd:2434:111  */
  assign n4840_o = n4839_o & n4836_o;
  /* TG68KdotC_Kernel.vhd:2435:104  */
  assign n4841_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2435:116  */
  assign n4843_o = n4841_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2435:94  */
  assign n4844_o = n4843_o & n4840_o;
  /* TG68KdotC_Kernel.vhd:2439:80  */
  assign n4845_o = exec[63];
  /* TG68KdotC_Kernel.vhd:2439:73  */
  assign n4847_o = n4845_o ? 7'b0000001 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2442:104  */
  assign n4849_o = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:2442:89  */
  assign n4850_o = n4849_o & nextpass;
  /* TG68KdotC_Kernel.vhd:2442:120  */
  assign n4851_o = opcode[6];
  /* TG68KdotC_Kernel.vhd:2442:123  */
  assign n4852_o = ~n4851_o;
  /* TG68KdotC_Kernel.vhd:2442:110  */
  assign n4853_o = n4852_o & n4850_o;
  /* TG68KdotC_Kernel.vhd:2442:73  */
  assign n4856_o = n4853_o ? 2'b11 : n2026_o;
  /* TG68KdotC_Kernel.vhd:2434:65  */
  assign n4858_o = n4894_o ? 1'b1 : n2015_o;
  assign n4859_o = n2162_o[1];
  assign n4860_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n4861_o = n2037_o ? n4859_o : n4860_o;
  /* TG68KdotC_Kernel.vhd:2442:73  */
  assign n4862_o = n4853_o ? 1'b1 : n4861_o;
  /* TG68KdotC_Kernel.vhd:2442:73  */
  assign n4864_o = n4853_o ? 7'b0011000 : n4847_o;
  /* TG68KdotC_Kernel.vhd:2449:87  */
  assign n4866_o = micro_state == 7'b0000101;
  /* TG68KdotC_Kernel.vhd:2449:106  */
  assign n4867_o = brief[8];
  /* TG68KdotC_Kernel.vhd:2449:109  */
  assign n4868_o = ~n4867_o;
  /* TG68KdotC_Kernel.vhd:2449:97  */
  assign n4869_o = n4868_o & n4866_o;
  /* TG68KdotC_Kernel.vhd:2449:73  */
  assign n4871_o = n4869_o ? 1'b1 : make_berr;
  /* TG68KdotC_Kernel.vhd:2452:81  */
  assign n4873_o = state == 2'b00;
  /* TG68KdotC_Kernel.vhd:2452:73  */
  assign n4876_o = n4873_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2456:79  */
  assign n4878_o = set[62];
  /* TG68KdotC_Kernel.vhd:2457:88  */
  assign n4879_o = exec[73];
  /* TG68KdotC_Kernel.vhd:2457:100  */
  assign n4880_o = ~n4879_o;
  /* TG68KdotC_Kernel.vhd:2457:105  */
  assign n4881_o = n4880_o | long_done;
  /* TG68KdotC_Kernel.vhd:2456:73  */
  assign n4883_o = n4885_o ? 1'b1 : n4871_o;
  /* TG68KdotC_Kernel.vhd:2456:73  */
  assign n4885_o = n4881_o & n4878_o;
  /* TG68KdotC_Kernel.vhd:2456:73  */
  assign n4887_o = n4878_o ? 2'b01 : n4856_o;
  assign n4888_o = n1909_o[63];
  /* TG68KdotC_Kernel.vhd:2456:73  */
  assign n4889_o = n4878_o ? 1'b1 : n4888_o;
  /* TG68KdotC_Kernel.vhd:2434:65  */
  assign n4890_o = n4844_o ? n4883_o : make_berr;
  /* TG68KdotC_Kernel.vhd:2434:65  */
  assign n4892_o = n4844_o ? 2'b10 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2434:65  */
  assign n4893_o = n4844_o ? n4887_o : n2026_o;
  /* TG68KdotC_Kernel.vhd:2434:65  */
  assign n4894_o = n4853_o & n4844_o;
  /* TG68KdotC_Kernel.vhd:2434:65  */
  assign n4896_o = n4844_o ? n4876_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2434:65  */
  assign n4899_o = n4844_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2434:65  */
  assign n4902_o = n4844_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2434:65  */
  assign n4905_o = n4844_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2434:65  */
  assign n4908_o = n4844_o ? 1'b1 : 1'b0;
  assign n4909_o = {1'b1, n4889_o};
  assign n4910_o = n2162_o[1];
  assign n4911_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n4912_o = n2037_o ? n4910_o : n4911_o;
  /* TG68KdotC_Kernel.vhd:2434:65  */
  assign n4913_o = n4844_o ? n4862_o : n4912_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n4914_o = n5462_o ? n4909_o : n2178_o;
  /* TG68KdotC_Kernel.vhd:2434:65  */
  assign n4915_o = n4844_o ? n4864_o : n2180_o;
  /* TG68KdotC_Kernel.vhd:2468:76  */
  assign n4916_o = opcode[6:0];
  /* TG68KdotC_Kernel.vhd:2469:73  */
  assign n4918_o = n4916_o == 7'b1000000;
  /* TG68KdotC_Kernel.vhd:2469:87  */
  assign n4920_o = n4916_o == 7'b1000001;
  /* TG68KdotC_Kernel.vhd:2469:87  */
  assign n4921_o = n4918_o | n4920_o;
  /* TG68KdotC_Kernel.vhd:2469:97  */
  assign n4923_o = n4916_o == 7'b1000010;
  /* TG68KdotC_Kernel.vhd:2469:97  */
  assign n4924_o = n4921_o | n4923_o;
  /* TG68KdotC_Kernel.vhd:2469:107  */
  assign n4926_o = n4916_o == 7'b1000011;
  /* TG68KdotC_Kernel.vhd:2469:107  */
  assign n4927_o = n4924_o | n4926_o;
  /* TG68KdotC_Kernel.vhd:2469:117  */
  assign n4929_o = n4916_o == 7'b1000100;
  /* TG68KdotC_Kernel.vhd:2469:117  */
  assign n4930_o = n4927_o | n4929_o;
  /* TG68KdotC_Kernel.vhd:2469:127  */
  assign n4932_o = n4916_o == 7'b1000101;
  /* TG68KdotC_Kernel.vhd:2469:127  */
  assign n4933_o = n4930_o | n4932_o;
  /* TG68KdotC_Kernel.vhd:2469:137  */
  assign n4935_o = n4916_o == 7'b1000110;
  /* TG68KdotC_Kernel.vhd:2469:137  */
  assign n4936_o = n4933_o | n4935_o;
  /* TG68KdotC_Kernel.vhd:2469:147  */
  assign n4938_o = n4916_o == 7'b1000111;
  /* TG68KdotC_Kernel.vhd:2469:147  */
  assign n4939_o = n4936_o | n4938_o;
  /* TG68KdotC_Kernel.vhd:2469:157  */
  assign n4941_o = n4916_o == 7'b1001000;
  /* TG68KdotC_Kernel.vhd:2469:157  */
  assign n4942_o = n4939_o | n4941_o;
  /* TG68KdotC_Kernel.vhd:2470:87  */
  assign n4944_o = n4916_o == 7'b1001001;
  /* TG68KdotC_Kernel.vhd:2470:87  */
  assign n4945_o = n4942_o | n4944_o;
  /* TG68KdotC_Kernel.vhd:2470:97  */
  assign n4947_o = n4916_o == 7'b1001010;
  /* TG68KdotC_Kernel.vhd:2470:97  */
  assign n4948_o = n4945_o | n4947_o;
  /* TG68KdotC_Kernel.vhd:2470:107  */
  assign n4950_o = n4916_o == 7'b1001011;
  /* TG68KdotC_Kernel.vhd:2470:107  */
  assign n4951_o = n4948_o | n4950_o;
  /* TG68KdotC_Kernel.vhd:2470:117  */
  assign n4953_o = n4916_o == 7'b1001100;
  /* TG68KdotC_Kernel.vhd:2470:117  */
  assign n4954_o = n4951_o | n4953_o;
  /* TG68KdotC_Kernel.vhd:2470:127  */
  assign n4956_o = n4916_o == 7'b1001101;
  /* TG68KdotC_Kernel.vhd:2470:127  */
  assign n4957_o = n4954_o | n4956_o;
  /* TG68KdotC_Kernel.vhd:2470:137  */
  assign n4959_o = n4916_o == 7'b1001110;
  /* TG68KdotC_Kernel.vhd:2470:137  */
  assign n4960_o = n4957_o | n4959_o;
  /* TG68KdotC_Kernel.vhd:2470:147  */
  assign n4962_o = n4916_o == 7'b1001111;
  /* TG68KdotC_Kernel.vhd:2470:147  */
  assign n4963_o = n4960_o | n4962_o;
  /* TG68KdotC_Kernel.vhd:2479:81  */
  assign n4971_o = decodeopc ? 1'b1 : n2015_o;
  /* TG68KdotC_Kernel.vhd:2479:81  */
  assign n4974_o = decodeopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2479:81  */
  assign n4977_o = decodeopc ? 1'b1 : 1'b0;
  assign n4978_o = n1909_o[44];
  /* TG68KdotC_Kernel.vhd:2479:81  */
  assign n4979_o = decodeopc ? 1'b1 : n4978_o;
  assign n4980_o = n2162_o[1];
  assign n4981_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n4982_o = n2037_o ? n4980_o : n4981_o;
  /* TG68KdotC_Kernel.vhd:2479:81  */
  assign n4983_o = decodeopc ? 1'b1 : n4982_o;
  assign n4984_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:2479:81  */
  assign n4985_o = decodeopc ? 1'b1 : n4984_o;
  /* TG68KdotC_Kernel.vhd:2479:81  */
  assign n4987_o = decodeopc ? 7'b0100011 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2474:73  */
  assign n4989_o = n4916_o == 7'b1010000;
  /* TG68KdotC_Kernel.vhd:2474:87  */
  assign n4991_o = n4916_o == 7'b1010001;
  /* TG68KdotC_Kernel.vhd:2474:87  */
  assign n4992_o = n4989_o | n4991_o;
  /* TG68KdotC_Kernel.vhd:2474:97  */
  assign n4994_o = n4916_o == 7'b1010010;
  /* TG68KdotC_Kernel.vhd:2474:97  */
  assign n4995_o = n4992_o | n4994_o;
  /* TG68KdotC_Kernel.vhd:2474:107  */
  assign n4997_o = n4916_o == 7'b1010011;
  /* TG68KdotC_Kernel.vhd:2474:107  */
  assign n4998_o = n4995_o | n4997_o;
  /* TG68KdotC_Kernel.vhd:2474:117  */
  assign n5000_o = n4916_o == 7'b1010100;
  /* TG68KdotC_Kernel.vhd:2474:117  */
  assign n5001_o = n4998_o | n5000_o;
  /* TG68KdotC_Kernel.vhd:2474:127  */
  assign n5003_o = n4916_o == 7'b1010101;
  /* TG68KdotC_Kernel.vhd:2474:127  */
  assign n5004_o = n5001_o | n5003_o;
  /* TG68KdotC_Kernel.vhd:2474:137  */
  assign n5006_o = n4916_o == 7'b1010110;
  /* TG68KdotC_Kernel.vhd:2474:137  */
  assign n5007_o = n5004_o | n5006_o;
  /* TG68KdotC_Kernel.vhd:2474:147  */
  assign n5009_o = n4916_o == 7'b1010111;
  /* TG68KdotC_Kernel.vhd:2474:147  */
  assign n5010_o = n5007_o | n5009_o;
  /* TG68KdotC_Kernel.vhd:2494:81  */
  assign n5017_o = decodeopc ? 2'b01 : n2026_o;
  /* TG68KdotC_Kernel.vhd:2494:81  */
  assign n5019_o = decodeopc ? 1'b1 : n2015_o;
  /* TG68KdotC_Kernel.vhd:2494:81  */
  assign n5022_o = decodeopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2494:81  */
  assign n5025_o = decodeopc ? 1'b1 : 1'b0;
  assign n5026_o = n1909_o[0];
  /* TG68KdotC_Kernel.vhd:2494:81  */
  assign n5027_o = decodeopc ? 1'b1 : n5026_o;
  assign n5028_o = n1909_o[34];
  /* TG68KdotC_Kernel.vhd:2494:81  */
  assign n5029_o = decodeopc ? 1'b1 : n5028_o;
  /* TG68KdotC_Kernel.vhd:2494:81  */
  assign n5031_o = decodeopc ? 7'b0100101 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2489:73  */
  assign n5033_o = n4916_o == 7'b1011000;
  /* TG68KdotC_Kernel.vhd:2489:87  */
  assign n5035_o = n4916_o == 7'b1011001;
  /* TG68KdotC_Kernel.vhd:2489:87  */
  assign n5036_o = n5033_o | n5035_o;
  /* TG68KdotC_Kernel.vhd:2489:97  */
  assign n5038_o = n4916_o == 7'b1011010;
  /* TG68KdotC_Kernel.vhd:2489:97  */
  assign n5039_o = n5036_o | n5038_o;
  /* TG68KdotC_Kernel.vhd:2489:107  */
  assign n5041_o = n4916_o == 7'b1011011;
  /* TG68KdotC_Kernel.vhd:2489:107  */
  assign n5042_o = n5039_o | n5041_o;
  /* TG68KdotC_Kernel.vhd:2489:117  */
  assign n5044_o = n4916_o == 7'b1011100;
  /* TG68KdotC_Kernel.vhd:2489:117  */
  assign n5045_o = n5042_o | n5044_o;
  /* TG68KdotC_Kernel.vhd:2489:127  */
  assign n5047_o = n4916_o == 7'b1011101;
  /* TG68KdotC_Kernel.vhd:2489:127  */
  assign n5048_o = n5045_o | n5047_o;
  /* TG68KdotC_Kernel.vhd:2489:137  */
  assign n5050_o = n4916_o == 7'b1011110;
  /* TG68KdotC_Kernel.vhd:2489:137  */
  assign n5051_o = n5048_o | n5050_o;
  /* TG68KdotC_Kernel.vhd:2489:147  */
  assign n5053_o = n4916_o == 7'b1011111;
  /* TG68KdotC_Kernel.vhd:2489:147  */
  assign n5054_o = n5051_o | n5053_o;
  /* TG68KdotC_Kernel.vhd:2505:81  */
  assign n5057_o = svmode ? 2'b10 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2505:81  */
  assign n5060_o = svmode ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2505:81  */
  assign n5063_o = svmode ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2505:81  */
  assign n5066_o = svmode ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2505:81  */
  assign n5069_o = svmode ? 1'b0 : 1'b1;
  assign n5070_o = n2017_o[0];
  assign n5071_o = n1909_o[65];
  /* TG68KdotC_Kernel.vhd:1578:17  */
  assign n5072_o = n2010_o ? n5070_o : n5071_o;
  /* TG68KdotC_Kernel.vhd:2505:81  */
  assign n5073_o = svmode ? 1'b1 : n5072_o;
  /* TG68KdotC_Kernel.vhd:2504:73  */
  assign n5075_o = n4916_o == 7'b1100000;
  /* TG68KdotC_Kernel.vhd:2504:87  */
  assign n5077_o = n4916_o == 7'b1100001;
  /* TG68KdotC_Kernel.vhd:2504:87  */
  assign n5078_o = n5075_o | n5077_o;
  /* TG68KdotC_Kernel.vhd:2504:97  */
  assign n5080_o = n4916_o == 7'b1100010;
  /* TG68KdotC_Kernel.vhd:2504:97  */
  assign n5081_o = n5078_o | n5080_o;
  /* TG68KdotC_Kernel.vhd:2504:107  */
  assign n5083_o = n4916_o == 7'b1100011;
  /* TG68KdotC_Kernel.vhd:2504:107  */
  assign n5084_o = n5081_o | n5083_o;
  /* TG68KdotC_Kernel.vhd:2504:117  */
  assign n5086_o = n4916_o == 7'b1100100;
  /* TG68KdotC_Kernel.vhd:2504:117  */
  assign n5087_o = n5084_o | n5086_o;
  /* TG68KdotC_Kernel.vhd:2504:127  */
  assign n5089_o = n4916_o == 7'b1100101;
  /* TG68KdotC_Kernel.vhd:2504:127  */
  assign n5090_o = n5087_o | n5089_o;
  /* TG68KdotC_Kernel.vhd:2504:137  */
  assign n5092_o = n4916_o == 7'b1100110;
  /* TG68KdotC_Kernel.vhd:2504:137  */
  assign n5093_o = n5090_o | n5092_o;
  /* TG68KdotC_Kernel.vhd:2504:147  */
  assign n5095_o = n4916_o == 7'b1100111;
  /* TG68KdotC_Kernel.vhd:2504:147  */
  assign n5096_o = n5093_o | n5095_o;
  /* TG68KdotC_Kernel.vhd:2517:81  */
  assign n5100_o = svmode ? 2'b10 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2517:81  */
  assign n5103_o = svmode ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2517:81  */
  assign n5106_o = svmode ? 1'b0 : 1'b1;
  assign n5107_o = n2017_o[1];
  assign n5108_o = n1909_o[66];
  /* TG68KdotC_Kernel.vhd:1578:17  */
  assign n5109_o = n2010_o ? n5107_o : n5108_o;
  /* TG68KdotC_Kernel.vhd:2517:81  */
  assign n5110_o = svmode ? 1'b1 : n5109_o;
  /* TG68KdotC_Kernel.vhd:2517:81  */
  assign n5112_o = svmode ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2516:73  */
  assign n5114_o = n4916_o == 7'b1101000;
  /* TG68KdotC_Kernel.vhd:2516:87  */
  assign n5116_o = n4916_o == 7'b1101001;
  /* TG68KdotC_Kernel.vhd:2516:87  */
  assign n5117_o = n5114_o | n5116_o;
  /* TG68KdotC_Kernel.vhd:2516:97  */
  assign n5119_o = n4916_o == 7'b1101010;
  /* TG68KdotC_Kernel.vhd:2516:97  */
  assign n5120_o = n5117_o | n5119_o;
  /* TG68KdotC_Kernel.vhd:2516:107  */
  assign n5122_o = n4916_o == 7'b1101011;
  /* TG68KdotC_Kernel.vhd:2516:107  */
  assign n5123_o = n5120_o | n5122_o;
  /* TG68KdotC_Kernel.vhd:2516:117  */
  assign n5125_o = n4916_o == 7'b1101100;
  /* TG68KdotC_Kernel.vhd:2516:117  */
  assign n5126_o = n5123_o | n5125_o;
  /* TG68KdotC_Kernel.vhd:2516:127  */
  assign n5128_o = n4916_o == 7'b1101101;
  /* TG68KdotC_Kernel.vhd:2516:127  */
  assign n5129_o = n5126_o | n5128_o;
  /* TG68KdotC_Kernel.vhd:2516:137  */
  assign n5131_o = n4916_o == 7'b1101110;
  /* TG68KdotC_Kernel.vhd:2516:137  */
  assign n5132_o = n5129_o | n5131_o;
  /* TG68KdotC_Kernel.vhd:2516:147  */
  assign n5134_o = n4916_o == 7'b1101111;
  /* TG68KdotC_Kernel.vhd:2516:147  */
  assign n5135_o = n5132_o | n5134_o;
  /* TG68KdotC_Kernel.vhd:2528:90  */
  assign n5136_o = ~svmode;
  /* TG68KdotC_Kernel.vhd:2533:89  */
  assign n5140_o = decodeopc ? 6'b000000 : n1906_o;
  assign n5141_o = n1909_o[24];
  /* TG68KdotC_Kernel.vhd:2533:89  */
  assign n5142_o = decodeopc ? 1'b1 : n5141_o;
  /* TG68KdotC_Kernel.vhd:2528:81  */
  assign n5143_o = n5136_o ? n1906_o : n5140_o;
  /* TG68KdotC_Kernel.vhd:2528:81  */
  assign n5146_o = n5136_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2528:81  */
  assign n5149_o = n5136_o ? 1'b1 : 1'b0;
  assign n5150_o = n1909_o[24];
  /* TG68KdotC_Kernel.vhd:2528:81  */
  assign n5151_o = n5136_o ? n5150_o : n5142_o;
  assign n5152_o = n1909_o[74];
  /* TG68KdotC_Kernel.vhd:2528:81  */
  assign n5153_o = n5136_o ? n5152_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:2527:73  */
  assign n5155_o = n4916_o == 7'b1110000;
  /* TG68KdotC_Kernel.vhd:2539:73  */
  assign n5157_o = n4916_o == 7'b1110001;
  /* TG68KdotC_Kernel.vhd:2542:90  */
  assign n5158_o = ~svmode;
  /* TG68KdotC_Kernel.vhd:2546:89  */
  assign n5160_o = decodeopc ? 1'b1 : n2148_o;
  /* TG68KdotC_Kernel.vhd:2546:89  */
  assign n5163_o = decodeopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2550:89  */
  assign n5165_o = stop ? 1'b1 : make_berr;
  /* TG68KdotC_Kernel.vhd:2542:81  */
  assign n5166_o = n5158_o ? make_berr : n5165_o;
  /* TG68KdotC_Kernel.vhd:2542:81  */
  assign n5167_o = n5158_o ? n2148_o : n5160_o;
  /* TG68KdotC_Kernel.vhd:2542:81  */
  assign n5170_o = n5158_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2542:81  */
  assign n5173_o = n5158_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2542:81  */
  assign n5175_o = n5158_o ? 1'b0 : n5163_o;
  /* TG68KdotC_Kernel.vhd:2541:73  */
  assign n5177_o = n4916_o == 7'b1110010;
  /* TG68KdotC_Kernel.vhd:2557:104  */
  assign n5178_o = opcode[2];
  /* TG68KdotC_Kernel.vhd:2557:95  */
  assign n5179_o = svmode | n5178_o;
  /* TG68KdotC_Kernel.vhd:2562:106  */
  assign n5181_o = opcode[2];
  assign n5184_o = n1909_o[59];
  /* TG68KdotC_Kernel.vhd:2562:97  */
  assign n5185_o = n5181_o ? n5184_o : 1'b1;
  assign n5186_o = n1909_o[60];
  /* TG68KdotC_Kernel.vhd:2562:97  */
  assign n5187_o = n5181_o ? 1'b1 : n5186_o;
  /* TG68KdotC_Kernel.vhd:2557:81  */
  assign n5189_o = n5201_o ? 2'b10 : n2026_o;
  /* TG68KdotC_Kernel.vhd:2557:81  */
  assign n5191_o = n5202_o ? 1'b1 : n2015_o;
  assign n5192_o = {n5187_o, n5185_o};
  assign n5193_o = n2162_o[0];
  assign n5194_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n5195_o = n2037_o ? n5193_o : n5194_o;
  /* TG68KdotC_Kernel.vhd:2558:89  */
  assign n5196_o = decodeopc ? 1'b1 : n5195_o;
  assign n5197_o = n1909_o[60:59];
  /* TG68KdotC_Kernel.vhd:2557:81  */
  assign n5198_o = n5214_o ? n5192_o : n5197_o;
  /* TG68KdotC_Kernel.vhd:2557:81  */
  assign n5200_o = n5215_o ? 7'b0101011 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2557:81  */
  assign n5201_o = decodeopc & n5179_o;
  /* TG68KdotC_Kernel.vhd:2557:81  */
  assign n5202_o = decodeopc & n5179_o;
  /* TG68KdotC_Kernel.vhd:2557:81  */
  assign n5205_o = n5179_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2557:81  */
  assign n5208_o = n5179_o ? 1'b0 : 1'b1;
  assign n5209_o = n2162_o[0];
  assign n5210_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n5211_o = n2037_o ? n5209_o : n5210_o;
  /* TG68KdotC_Kernel.vhd:2557:81  */
  assign n5212_o = n5179_o ? n5196_o : n5211_o;
  /* TG68KdotC_Kernel.vhd:2557:81  */
  assign n5214_o = decodeopc & n5179_o;
  /* TG68KdotC_Kernel.vhd:2557:81  */
  assign n5215_o = decodeopc & n5179_o;
  /* TG68KdotC_Kernel.vhd:2556:73  */
  assign n5217_o = n4916_o == 7'b1110011;
  /* TG68KdotC_Kernel.vhd:2556:87  */
  assign n5219_o = n4916_o == 7'b1110111;
  /* TG68KdotC_Kernel.vhd:2556:87  */
  assign n5220_o = n5217_o | n5219_o;
  /* TG68KdotC_Kernel.vhd:2576:81  */
  assign n5225_o = decodeopc ? 2'b10 : n2026_o;
  /* TG68KdotC_Kernel.vhd:2576:81  */
  assign n5227_o = decodeopc ? 1'b1 : n2015_o;
  /* TG68KdotC_Kernel.vhd:2576:81  */
  assign n5229_o = decodeopc ? 1'b1 : n2154_o;
  assign n5230_o = {1'b1, 1'b1};
  assign n5231_o = n2162_o[0];
  assign n5232_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n5233_o = n2037_o ? n5231_o : n5232_o;
  /* TG68KdotC_Kernel.vhd:2576:81  */
  assign n5234_o = decodeopc ? 1'b1 : n5233_o;
  assign n5235_o = n1909_o[58:57];
  /* TG68KdotC_Kernel.vhd:2576:81  */
  assign n5236_o = decodeopc ? n5230_o : n5235_o;
  /* TG68KdotC_Kernel.vhd:2576:81  */
  assign n5238_o = decodeopc ? 7'b0110000 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2574:73  */
  assign n5240_o = n4916_o == 7'b1110100;
  /* TG68KdotC_Kernel.vhd:2589:81  */
  assign n5245_o = decodeopc ? 2'b10 : n2026_o;
  /* TG68KdotC_Kernel.vhd:2589:81  */
  assign n5247_o = decodeopc ? 1'b1 : n2015_o;
  assign n5248_o = {1'b1, 1'b1};
  assign n5249_o = n2162_o[0];
  assign n5250_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n5251_o = n2037_o ? n5249_o : n5250_o;
  /* TG68KdotC_Kernel.vhd:2589:81  */
  assign n5252_o = decodeopc ? 1'b1 : n5251_o;
  assign n5253_o = n1909_o[58:57];
  /* TG68KdotC_Kernel.vhd:2589:81  */
  assign n5254_o = decodeopc ? n5248_o : n5253_o;
  /* TG68KdotC_Kernel.vhd:2589:81  */
  assign n5256_o = decodeopc ? 7'b0011000 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2587:73  */
  assign n5258_o = n4916_o == 7'b1110101;
  /* TG68KdotC_Kernel.vhd:2599:81  */
  assign n5260_o = decodeopc ? 2'b01 : n2026_o;
  /* TG68KdotC_Kernel.vhd:2602:89  */
  assign n5261_o = flags[1];
  /* TG68KdotC_Kernel.vhd:2602:106  */
  assign n5263_o = state == 2'b01;
  /* TG68KdotC_Kernel.vhd:2602:97  */
  assign n5264_o = n5263_o & n5261_o;
  /* TG68KdotC_Kernel.vhd:2602:81  */
  assign n5267_o = n5264_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2602:81  */
  assign n5270_o = n5264_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2598:73  */
  assign n5272_o = n4916_o == 7'b1110110;
  /* TG68KdotC_Kernel.vhd:2608:87  */
  assign n5274_o = cpu == 2'b00;
  /* TG68KdotC_Kernel.vhd:2611:93  */
  assign n5275_o = ~svmode;
  /* TG68KdotC_Kernel.vhd:2616:106  */
  assign n5276_o = last_data_read[11:0];
  /* TG68KdotC_Kernel.vhd:2616:119  */
  assign n5278_o = n5276_o == 12'b100000000000;
  /* TG68KdotC_Kernel.vhd:2618:106  */
  assign n5280_o = opcode[0];
  assign n5282_o = n2017_o[0];
  assign n5283_o = n1909_o[65];
  /* TG68KdotC_Kernel.vhd:1578:17  */
  assign n5284_o = n2010_o ? n5282_o : n5283_o;
  /* TG68KdotC_Kernel.vhd:2618:97  */
  assign n5285_o = n5280_o ? 1'b1 : n5284_o;
  assign n5286_o = {1'b1, n5285_o};
  /* TG68KdotC_Kernel.vhd:2616:89  */
  assign n5287_o = n5278_o ? n5286_o : n2019_o;
  /* TG68KdotC_Kernel.vhd:2622:98  */
  assign n5288_o = opcode[0];
  /* TG68KdotC_Kernel.vhd:2622:101  */
  assign n5289_o = ~n5288_o;
  /* TG68KdotC_Kernel.vhd:2622:89  */
  assign n5293_o = n5289_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2622:89  */
  assign n5295_o = n5289_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2627:89  */
  assign n5297_o = decodeopc ? 1'b1 : n2151_o;
  /* TG68KdotC_Kernel.vhd:2627:89  */
  assign n5299_o = decodeopc ? 7'b1001101 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2611:81  */
  assign n5301_o = n5275_o ? n1921_o : 2'b10;
  /* TG68KdotC_Kernel.vhd:2611:81  */
  assign n5302_o = n5275_o ? n2151_o : n5297_o;
  /* TG68KdotC_Kernel.vhd:2611:81  */
  assign n5305_o = n5275_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2611:81  */
  assign n5308_o = n5275_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2611:81  */
  assign n5309_o = n5275_o ? n2019_o : n5287_o;
  assign n5310_o = {n5295_o, n5293_o};
  /* TG68KdotC_Kernel.vhd:2611:81  */
  assign n5312_o = n5275_o ? 2'b00 : n5310_o;
  /* TG68KdotC_Kernel.vhd:2611:81  */
  assign n5313_o = n5275_o ? n2180_o : n5299_o;
  /* TG68KdotC_Kernel.vhd:2608:81  */
  assign n5314_o = n5274_o ? n1921_o : n5301_o;
  /* TG68KdotC_Kernel.vhd:2608:81  */
  assign n5315_o = n5274_o ? n2151_o : n5302_o;
  /* TG68KdotC_Kernel.vhd:2608:81  */
  assign n5318_o = n5274_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2608:81  */
  assign n5320_o = n5274_o ? 1'b0 : n5305_o;
  /* TG68KdotC_Kernel.vhd:2608:81  */
  assign n5322_o = n5274_o ? 1'b1 : n5308_o;
  /* TG68KdotC_Kernel.vhd:2608:81  */
  assign n5323_o = n5274_o ? n2019_o : n5309_o;
  /* TG68KdotC_Kernel.vhd:2608:81  */
  assign n5325_o = n5274_o ? 2'b00 : n5312_o;
  /* TG68KdotC_Kernel.vhd:2608:81  */
  assign n5326_o = n5274_o ? n2180_o : n5313_o;
  /* TG68KdotC_Kernel.vhd:2607:73  */
  assign n5328_o = n4916_o == 7'b1111010;
  /* TG68KdotC_Kernel.vhd:2607:87  */
  assign n5330_o = n4916_o == 7'b1111011;
  /* TG68KdotC_Kernel.vhd:2607:87  */
  assign n5331_o = n5328_o | n5330_o;
  assign n5332_o = {n5331_o, n5272_o, n5258_o, n5240_o, n5220_o, n5177_o, n5157_o, n5155_o, n5135_o, n5096_o, n5054_o, n5010_o, n4963_o};
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5333_o = make_berr;
      13'b0100000000000: n5333_o = make_berr;
      13'b0010000000000: n5333_o = make_berr;
      13'b0001000000000: n5333_o = make_berr;
      13'b0000100000000: n5333_o = make_berr;
      13'b0000010000000: n5333_o = n5166_o;
      13'b0000001000000: n5333_o = make_berr;
      13'b0000000100000: n5333_o = make_berr;
      13'b0000000010000: n5333_o = make_berr;
      13'b0000000001000: n5333_o = make_berr;
      13'b0000000000100: n5333_o = make_berr;
      13'b0000000000010: n5333_o = make_berr;
      13'b0000000000001: n5333_o = make_berr;
      default: n5333_o = make_berr;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5338_o = n5314_o;
      13'b0100000000000: n5338_o = n1921_o;
      13'b0010000000000: n5338_o = 2'b10;
      13'b0001000000000: n5338_o = 2'b10;
      13'b0000100000000: n5338_o = n1921_o;
      13'b0000010000000: n5338_o = n1921_o;
      13'b0000001000000: n5338_o = n1921_o;
      13'b0000000100000: n5338_o = n1921_o;
      13'b0000000010000: n5338_o = n5100_o;
      13'b0000000001000: n5338_o = n5057_o;
      13'b0000000000100: n5338_o = 2'b10;
      13'b0000000000010: n5338_o = 2'b10;
      13'b0000000000001: n5338_o = n1921_o;
      default: n5338_o = n1921_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5339_o = n2026_o;
      13'b0100000000000: n5339_o = n5260_o;
      13'b0010000000000: n5339_o = n5245_o;
      13'b0001000000000: n5339_o = n5225_o;
      13'b0000100000000: n5339_o = n5189_o;
      13'b0000010000000: n5339_o = n2026_o;
      13'b0000001000000: n5339_o = n2026_o;
      13'b0000000100000: n5339_o = n2026_o;
      13'b0000000010000: n5339_o = n2026_o;
      13'b0000000001000: n5339_o = n2026_o;
      13'b0000000000100: n5339_o = n5017_o;
      13'b0000000000010: n5339_o = n2026_o;
      13'b0000000000001: n5339_o = n2026_o;
      default: n5339_o = n2026_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5340_o = n2148_o;
      13'b0100000000000: n5340_o = n2148_o;
      13'b0010000000000: n5340_o = n2148_o;
      13'b0001000000000: n5340_o = n2148_o;
      13'b0000100000000: n5340_o = n2148_o;
      13'b0000010000000: n5340_o = n5167_o;
      13'b0000001000000: n5340_o = n2148_o;
      13'b0000000100000: n5340_o = n2148_o;
      13'b0000000010000: n5340_o = n2148_o;
      13'b0000000001000: n5340_o = n2148_o;
      13'b0000000000100: n5340_o = n2148_o;
      13'b0000000000010: n5340_o = n2148_o;
      13'b0000000000001: n5340_o = n2148_o;
      default: n5340_o = n2148_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5341_o = n5315_o;
      13'b0100000000000: n5341_o = n2151_o;
      13'b0010000000000: n5341_o = n2151_o;
      13'b0001000000000: n5341_o = n2151_o;
      13'b0000100000000: n5341_o = n2151_o;
      13'b0000010000000: n5341_o = n2151_o;
      13'b0000001000000: n5341_o = n2151_o;
      13'b0000000100000: n5341_o = n2151_o;
      13'b0000000010000: n5341_o = n2151_o;
      13'b0000000001000: n5341_o = n2151_o;
      13'b0000000000100: n5341_o = n2151_o;
      13'b0000000000010: n5341_o = n2151_o;
      13'b0000000000001: n5341_o = n2151_o;
      default: n5341_o = n2151_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5342_o = n2015_o;
      13'b0100000000000: n5342_o = n2015_o;
      13'b0010000000000: n5342_o = n5247_o;
      13'b0001000000000: n5342_o = n5227_o;
      13'b0000100000000: n5342_o = n5191_o;
      13'b0000010000000: n5342_o = n2015_o;
      13'b0000001000000: n5342_o = n2015_o;
      13'b0000000100000: n5342_o = n2015_o;
      13'b0000000010000: n5342_o = n2015_o;
      13'b0000000001000: n5342_o = n2015_o;
      13'b0000000000100: n5342_o = n5019_o;
      13'b0000000000010: n5342_o = n4971_o;
      13'b0000000000001: n5342_o = n2015_o;
      default: n5342_o = n2015_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5344_o = 1'b0;
      13'b0100000000000: n5344_o = 1'b0;
      13'b0010000000000: n5344_o = 1'b0;
      13'b0001000000000: n5344_o = 1'b0;
      13'b0000100000000: n5344_o = 1'b0;
      13'b0000010000000: n5344_o = 1'b0;
      13'b0000001000000: n5344_o = 1'b0;
      13'b0000000100000: n5344_o = 1'b0;
      13'b0000000010000: n5344_o = 1'b0;
      13'b0000000001000: n5344_o = n5060_o;
      13'b0000000000100: n5344_o = n5022_o;
      13'b0000000000010: n5344_o = n4974_o;
      13'b0000000000001: n5344_o = 1'b0;
      default: n5344_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5346_o = 1'b0;
      13'b0100000000000: n5346_o = 1'b0;
      13'b0010000000000: n5346_o = 1'b0;
      13'b0001000000000: n5346_o = 1'b0;
      13'b0000100000000: n5346_o = 1'b0;
      13'b0000010000000: n5346_o = 1'b0;
      13'b0000001000000: n5346_o = 1'b0;
      13'b0000000100000: n5346_o = 1'b0;
      13'b0000000010000: n5346_o = 1'b0;
      13'b0000000001000: n5346_o = n5063_o;
      13'b0000000000100: n5346_o = n5025_o;
      13'b0000000000010: n5346_o = n4977_o;
      13'b0000000000001: n5346_o = 1'b0;
      default: n5346_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5347_o = n1906_o;
      13'b0100000000000: n5347_o = n1906_o;
      13'b0010000000000: n5347_o = n1906_o;
      13'b0001000000000: n5347_o = n1906_o;
      13'b0000100000000: n5347_o = n1906_o;
      13'b0000010000000: n5347_o = n1906_o;
      13'b0000001000000: n5347_o = n1906_o;
      13'b0000000100000: n5347_o = n5143_o;
      13'b0000000010000: n5347_o = n1906_o;
      13'b0000000001000: n5347_o = n1906_o;
      13'b0000000000100: n5347_o = n1906_o;
      13'b0000000000010: n5347_o = n1906_o;
      13'b0000000000001: n5347_o = n1906_o;
      default: n5347_o = n1906_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5348_o = n2154_o;
      13'b0100000000000: n5348_o = n2154_o;
      13'b0010000000000: n5348_o = n2154_o;
      13'b0001000000000: n5348_o = n5229_o;
      13'b0000100000000: n5348_o = n2154_o;
      13'b0000010000000: n5348_o = n2154_o;
      13'b0000001000000: n5348_o = n2154_o;
      13'b0000000100000: n5348_o = n2154_o;
      13'b0000000010000: n5348_o = n2154_o;
      13'b0000000001000: n5348_o = n2154_o;
      13'b0000000000100: n5348_o = n2154_o;
      13'b0000000000010: n5348_o = n2154_o;
      13'b0000000000001: n5348_o = n2154_o;
      default: n5348_o = n2154_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5351_o = n5318_o;
      13'b0100000000000: n5351_o = 1'b0;
      13'b0010000000000: n5351_o = 1'b0;
      13'b0001000000000: n5351_o = 1'b0;
      13'b0000100000000: n5351_o = 1'b0;
      13'b0000010000000: n5351_o = 1'b0;
      13'b0000001000000: n5351_o = 1'b0;
      13'b0000000100000: n5351_o = 1'b0;
      13'b0000000010000: n5351_o = 1'b0;
      13'b0000000001000: n5351_o = 1'b0;
      13'b0000000000100: n5351_o = 1'b0;
      13'b0000000000010: n5351_o = 1'b0;
      13'b0000000000001: n5351_o = 1'b0;
      default: n5351_o = 1'b1;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5353_o = n5320_o;
      13'b0100000000000: n5353_o = 1'b0;
      13'b0010000000000: n5353_o = 1'b0;
      13'b0001000000000: n5353_o = 1'b0;
      13'b0000100000000: n5353_o = n5205_o;
      13'b0000010000000: n5353_o = n5170_o;
      13'b0000001000000: n5353_o = 1'b0;
      13'b0000000100000: n5353_o = n5146_o;
      13'b0000000010000: n5353_o = n5103_o;
      13'b0000000001000: n5353_o = n5066_o;
      13'b0000000000100: n5353_o = 1'b0;
      13'b0000000000010: n5353_o = 1'b0;
      13'b0000000000001: n5353_o = 1'b0;
      default: n5353_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5356_o = 1'b0;
      13'b0100000000000: n5356_o = 1'b0;
      13'b0010000000000: n5356_o = 1'b0;
      13'b0001000000000: n5356_o = 1'b0;
      13'b0000100000000: n5356_o = 1'b0;
      13'b0000010000000: n5356_o = 1'b0;
      13'b0000001000000: n5356_o = 1'b0;
      13'b0000000100000: n5356_o = 1'b0;
      13'b0000000010000: n5356_o = 1'b0;
      13'b0000000001000: n5356_o = 1'b0;
      13'b0000000000100: n5356_o = 1'b0;
      13'b0000000000010: n5356_o = 1'b0;
      13'b0000000000001: n5356_o = 1'b1;
      default: n5356_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5358_o = 1'b0;
      13'b0100000000000: n5358_o = n5267_o;
      13'b0010000000000: n5358_o = 1'b0;
      13'b0001000000000: n5358_o = 1'b0;
      13'b0000100000000: n5358_o = 1'b0;
      13'b0000010000000: n5358_o = 1'b0;
      13'b0000001000000: n5358_o = 1'b0;
      13'b0000000100000: n5358_o = 1'b0;
      13'b0000000010000: n5358_o = 1'b0;
      13'b0000000001000: n5358_o = 1'b0;
      13'b0000000000100: n5358_o = 1'b0;
      13'b0000000000010: n5358_o = 1'b0;
      13'b0000000000001: n5358_o = 1'b0;
      default: n5358_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5362_o = n5322_o;
      13'b0100000000000: n5362_o = n5270_o;
      13'b0010000000000: n5362_o = 1'b0;
      13'b0001000000000: n5362_o = 1'b0;
      13'b0000100000000: n5362_o = n5208_o;
      13'b0000010000000: n5362_o = n5173_o;
      13'b0000001000000: n5362_o = 1'b0;
      13'b0000000100000: n5362_o = n5149_o;
      13'b0000000010000: n5362_o = n5106_o;
      13'b0000000001000: n5362_o = n5069_o;
      13'b0000000000100: n5362_o = 1'b0;
      13'b0000000000010: n5362_o = 1'b0;
      13'b0000000000001: n5362_o = 1'b1;
      default: n5362_o = 1'b1;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5364_o = 1'b0;
      13'b0100000000000: n5364_o = 1'b0;
      13'b0010000000000: n5364_o = 1'b0;
      13'b0001000000000: n5364_o = 1'b0;
      13'b0000100000000: n5364_o = 1'b0;
      13'b0000010000000: n5364_o = n5175_o;
      13'b0000001000000: n5364_o = 1'b0;
      13'b0000000100000: n5364_o = 1'b0;
      13'b0000000010000: n5364_o = 1'b0;
      13'b0000000001000: n5364_o = 1'b0;
      13'b0000000000100: n5364_o = 1'b0;
      13'b0000000000010: n5364_o = 1'b0;
      13'b0000000000001: n5364_o = 1'b0;
      default: n5364_o = 1'b0;
    endcase
  assign n5365_o = n1909_o[0];
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5366_o = n5365_o;
      13'b0100000000000: n5366_o = n5365_o;
      13'b0010000000000: n5366_o = n5365_o;
      13'b0001000000000: n5366_o = n5365_o;
      13'b0000100000000: n5366_o = n5365_o;
      13'b0000010000000: n5366_o = n5365_o;
      13'b0000001000000: n5366_o = n5365_o;
      13'b0000000100000: n5366_o = n5365_o;
      13'b0000000010000: n5366_o = n5365_o;
      13'b0000000001000: n5366_o = n5365_o;
      13'b0000000000100: n5366_o = n5027_o;
      13'b0000000000010: n5366_o = n5365_o;
      13'b0000000000001: n5366_o = n5365_o;
      default: n5366_o = n5365_o;
    endcase
  assign n5367_o = n1909_o[24];
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5368_o = n5367_o;
      13'b0100000000000: n5368_o = n5367_o;
      13'b0010000000000: n5368_o = n5367_o;
      13'b0001000000000: n5368_o = n5367_o;
      13'b0000100000000: n5368_o = n5367_o;
      13'b0000010000000: n5368_o = n5367_o;
      13'b0000001000000: n5368_o = n5367_o;
      13'b0000000100000: n5368_o = n5151_o;
      13'b0000000010000: n5368_o = n5367_o;
      13'b0000000001000: n5368_o = n5367_o;
      13'b0000000000100: n5368_o = n5367_o;
      13'b0000000000010: n5368_o = n5367_o;
      13'b0000000000001: n5368_o = n5367_o;
      default: n5368_o = n5367_o;
    endcase
  assign n5369_o = n1909_o[34];
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5370_o = n5369_o;
      13'b0100000000000: n5370_o = n5369_o;
      13'b0010000000000: n5370_o = n5369_o;
      13'b0001000000000: n5370_o = n5369_o;
      13'b0000100000000: n5370_o = n5369_o;
      13'b0000010000000: n5370_o = n5369_o;
      13'b0000001000000: n5370_o = n5369_o;
      13'b0000000100000: n5370_o = n5369_o;
      13'b0000000010000: n5370_o = n5369_o;
      13'b0000000001000: n5370_o = n5369_o;
      13'b0000000000100: n5370_o = n5029_o;
      13'b0000000000010: n5370_o = n5369_o;
      13'b0000000000001: n5370_o = n5369_o;
      default: n5370_o = n5369_o;
    endcase
  assign n5371_o = n1909_o[44];
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5372_o = n5371_o;
      13'b0100000000000: n5372_o = n5371_o;
      13'b0010000000000: n5372_o = n5371_o;
      13'b0001000000000: n5372_o = n5371_o;
      13'b0000100000000: n5372_o = n5371_o;
      13'b0000010000000: n5372_o = n5371_o;
      13'b0000001000000: n5372_o = n5371_o;
      13'b0000000100000: n5372_o = n5371_o;
      13'b0000000010000: n5372_o = n5371_o;
      13'b0000000001000: n5372_o = n5371_o;
      13'b0000000000100: n5372_o = n5371_o;
      13'b0000000000010: n5372_o = n4979_o;
      13'b0000000000001: n5372_o = n5371_o;
      default: n5372_o = n5371_o;
    endcase
  assign n5373_o = n2162_o[0];
  assign n5374_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n5375_o = n2037_o ? n5373_o : n5374_o;
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5376_o = n5375_o;
      13'b0100000000000: n5376_o = n5375_o;
      13'b0010000000000: n5376_o = n5252_o;
      13'b0001000000000: n5376_o = n5234_o;
      13'b0000100000000: n5376_o = n5212_o;
      13'b0000010000000: n5376_o = n5375_o;
      13'b0000001000000: n5376_o = n5375_o;
      13'b0000000100000: n5376_o = n5375_o;
      13'b0000000010000: n5376_o = n5375_o;
      13'b0000000001000: n5376_o = n5375_o;
      13'b0000000000100: n5376_o = n5375_o;
      13'b0000000000010: n5376_o = n5375_o;
      13'b0000000000001: n5376_o = n5375_o;
      default: n5376_o = n5375_o;
    endcase
  assign n5377_o = n2162_o[1];
  assign n5378_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n5379_o = n2037_o ? n5377_o : n5378_o;
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5380_o = n5379_o;
      13'b0100000000000: n5380_o = n5379_o;
      13'b0010000000000: n5380_o = n5379_o;
      13'b0001000000000: n5380_o = n5379_o;
      13'b0000100000000: n5380_o = n5379_o;
      13'b0000010000000: n5380_o = n5379_o;
      13'b0000001000000: n5380_o = n5379_o;
      13'b0000000100000: n5380_o = n5379_o;
      13'b0000000010000: n5380_o = n5379_o;
      13'b0000000001000: n5380_o = n5379_o;
      13'b0000000000100: n5380_o = n5379_o;
      13'b0000000000010: n5380_o = n4983_o;
      13'b0000000000001: n5380_o = n5379_o;
      default: n5380_o = n5379_o;
    endcase
  assign n5381_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5382_o = n5381_o;
      13'b0100000000000: n5382_o = n5381_o;
      13'b0010000000000: n5382_o = n5381_o;
      13'b0001000000000: n5382_o = n5381_o;
      13'b0000100000000: n5382_o = n5381_o;
      13'b0000010000000: n5382_o = n5381_o;
      13'b0000001000000: n5382_o = n5381_o;
      13'b0000000100000: n5382_o = n5381_o;
      13'b0000000010000: n5382_o = n5381_o;
      13'b0000000001000: n5382_o = n5381_o;
      13'b0000000000100: n5382_o = 1'b1;
      13'b0000000000010: n5382_o = 1'b1;
      13'b0000000000001: n5382_o = n5381_o;
      default: n5382_o = n5381_o;
    endcase
  assign n5383_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5384_o = n5383_o;
      13'b0100000000000: n5384_o = n5383_o;
      13'b0010000000000: n5384_o = n5383_o;
      13'b0001000000000: n5384_o = n5383_o;
      13'b0000100000000: n5384_o = n5383_o;
      13'b0000010000000: n5384_o = n5383_o;
      13'b0000001000000: n5384_o = n5383_o;
      13'b0000000100000: n5384_o = n5383_o;
      13'b0000000010000: n5384_o = n5383_o;
      13'b0000000001000: n5384_o = n5383_o;
      13'b0000000000100: n5384_o = n5383_o;
      13'b0000000000010: n5384_o = n4985_o;
      13'b0000000000001: n5384_o = n5383_o;
      default: n5384_o = n5383_o;
    endcase
  assign n5385_o = n1909_o[58:57];
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5386_o = n5385_o;
      13'b0100000000000: n5386_o = n5385_o;
      13'b0010000000000: n5386_o = n5254_o;
      13'b0001000000000: n5386_o = n5236_o;
      13'b0000100000000: n5386_o = n5385_o;
      13'b0000010000000: n5386_o = n5385_o;
      13'b0000001000000: n5386_o = n5385_o;
      13'b0000000100000: n5386_o = n5385_o;
      13'b0000000010000: n5386_o = n5385_o;
      13'b0000000001000: n5386_o = n5385_o;
      13'b0000000000100: n5386_o = n5385_o;
      13'b0000000000010: n5386_o = n5385_o;
      13'b0000000000001: n5386_o = n5385_o;
      default: n5386_o = n5385_o;
    endcase
  assign n5387_o = n1909_o[60:59];
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5388_o = n5387_o;
      13'b0100000000000: n5388_o = n5387_o;
      13'b0010000000000: n5388_o = n5387_o;
      13'b0001000000000: n5388_o = n5387_o;
      13'b0000100000000: n5388_o = n5198_o;
      13'b0000010000000: n5388_o = n5387_o;
      13'b0000001000000: n5388_o = n5387_o;
      13'b0000000100000: n5388_o = n5387_o;
      13'b0000000010000: n5388_o = n5387_o;
      13'b0000000001000: n5388_o = n5387_o;
      13'b0000000000100: n5388_o = n5387_o;
      13'b0000000000010: n5388_o = n5387_o;
      13'b0000000000001: n5388_o = n5387_o;
      default: n5388_o = n5387_o;
    endcase
  assign n5389_o = n5323_o[0];
  assign n5390_o = n2017_o[0];
  assign n5391_o = n1909_o[65];
  /* TG68KdotC_Kernel.vhd:1578:17  */
  assign n5392_o = n2010_o ? n5390_o : n5391_o;
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5393_o = n5389_o;
      13'b0100000000000: n5393_o = n5392_o;
      13'b0010000000000: n5393_o = n5392_o;
      13'b0001000000000: n5393_o = n5392_o;
      13'b0000100000000: n5393_o = n5392_o;
      13'b0000010000000: n5393_o = n5392_o;
      13'b0000001000000: n5393_o = n5392_o;
      13'b0000000100000: n5393_o = n5392_o;
      13'b0000000010000: n5393_o = n5392_o;
      13'b0000000001000: n5393_o = n5073_o;
      13'b0000000000100: n5393_o = n5392_o;
      13'b0000000000010: n5393_o = n5392_o;
      13'b0000000000001: n5393_o = n5392_o;
      default: n5393_o = n5392_o;
    endcase
  assign n5394_o = n5323_o[1];
  assign n5395_o = n2017_o[1];
  assign n5396_o = n1909_o[66];
  /* TG68KdotC_Kernel.vhd:1578:17  */
  assign n5397_o = n2010_o ? n5395_o : n5396_o;
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5398_o = n5394_o;
      13'b0100000000000: n5398_o = n5397_o;
      13'b0010000000000: n5398_o = n5397_o;
      13'b0001000000000: n5398_o = n5397_o;
      13'b0000100000000: n5398_o = n5397_o;
      13'b0000010000000: n5398_o = n5397_o;
      13'b0000001000000: n5398_o = n5397_o;
      13'b0000000100000: n5398_o = n5397_o;
      13'b0000000010000: n5398_o = n5110_o;
      13'b0000000001000: n5398_o = n5397_o;
      13'b0000000000100: n5398_o = n5397_o;
      13'b0000000000010: n5398_o = n5397_o;
      13'b0000000000001: n5398_o = n5397_o;
      default: n5398_o = n5397_o;
    endcase
  assign n5399_o = n1909_o[74];
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5400_o = n5399_o;
      13'b0100000000000: n5400_o = n5399_o;
      13'b0010000000000: n5400_o = n5399_o;
      13'b0001000000000: n5400_o = n5399_o;
      13'b0000100000000: n5400_o = n5399_o;
      13'b0000010000000: n5400_o = n5399_o;
      13'b0000001000000: n5400_o = n5399_o;
      13'b0000000100000: n5400_o = n5153_o;
      13'b0000000010000: n5400_o = n5399_o;
      13'b0000000001000: n5400_o = n5399_o;
      13'b0000000000100: n5400_o = n5399_o;
      13'b0000000000010: n5400_o = n5399_o;
      13'b0000000000001: n5400_o = n5399_o;
      default: n5400_o = n5399_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5402_o = 1'b0;
      13'b0100000000000: n5402_o = 1'b0;
      13'b0010000000000: n5402_o = 1'b0;
      13'b0001000000000: n5402_o = 1'b0;
      13'b0000100000000: n5402_o = 1'b0;
      13'b0000010000000: n5402_o = 1'b0;
      13'b0000001000000: n5402_o = 1'b0;
      13'b0000000100000: n5402_o = 1'b0;
      13'b0000000010000: n5402_o = 1'b0;
      13'b0000000001000: n5402_o = 1'b0;
      13'b0000000000100: n5402_o = 1'b1;
      13'b0000000000010: n5402_o = 1'b0;
      13'b0000000000001: n5402_o = 1'b0;
      default: n5402_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5404_o = 1'b0;
      13'b0100000000000: n5404_o = 1'b0;
      13'b0010000000000: n5404_o = 1'b0;
      13'b0001000000000: n5404_o = 1'b0;
      13'b0000100000000: n5404_o = 1'b0;
      13'b0000010000000: n5404_o = 1'b0;
      13'b0000001000000: n5404_o = 1'b0;
      13'b0000000100000: n5404_o = 1'b0;
      13'b0000000010000: n5404_o = 1'b0;
      13'b0000000001000: n5404_o = 1'b0;
      13'b0000000000100: n5404_o = 1'b0;
      13'b0000000000010: n5404_o = 1'b1;
      13'b0000000000001: n5404_o = 1'b0;
      default: n5404_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5406_o = n5325_o;
      13'b0100000000000: n5406_o = 2'b00;
      13'b0010000000000: n5406_o = 2'b00;
      13'b0001000000000: n5406_o = 2'b00;
      13'b0000100000000: n5406_o = 2'b00;
      13'b0000010000000: n5406_o = 2'b00;
      13'b0000001000000: n5406_o = 2'b00;
      13'b0000000100000: n5406_o = 2'b00;
      13'b0000000010000: n5406_o = 2'b00;
      13'b0000000001000: n5406_o = 2'b00;
      13'b0000000000100: n5406_o = 2'b00;
      13'b0000000000010: n5406_o = 2'b00;
      13'b0000000000001: n5406_o = 2'b00;
      default: n5406_o = 2'b00;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5408_o = 1'b0;
      13'b0100000000000: n5408_o = 1'b0;
      13'b0010000000000: n5408_o = 1'b0;
      13'b0001000000000: n5408_o = 1'b0;
      13'b0000100000000: n5408_o = 1'b0;
      13'b0000010000000: n5408_o = 1'b0;
      13'b0000001000000: n5408_o = 1'b0;
      13'b0000000100000: n5408_o = 1'b0;
      13'b0000000010000: n5408_o = n5112_o;
      13'b0000000001000: n5408_o = 1'b0;
      13'b0000000000100: n5408_o = 1'b1;
      13'b0000000000010: n5408_o = 1'b1;
      13'b0000000000001: n5408_o = 1'b0;
      default: n5408_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2468:65  */
  always @*
    case (n5332_o)
      13'b1000000000000: n5409_o = n5326_o;
      13'b0100000000000: n5409_o = n2180_o;
      13'b0010000000000: n5409_o = n5256_o;
      13'b0001000000000: n5409_o = n5238_o;
      13'b0000100000000: n5409_o = n5200_o;
      13'b0000010000000: n5409_o = n2180_o;
      13'b0000001000000: n5409_o = n2180_o;
      13'b0000000100000: n5409_o = n2180_o;
      13'b0000000010000: n5409_o = n2180_o;
      13'b0000000001000: n5409_o = n2180_o;
      13'b0000000000100: n5409_o = n5031_o;
      13'b0000000000010: n5409_o = n4987_o;
      13'b0000000000001: n5409_o = n2180_o;
      default: n5409_o = n2180_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5410_o = n4831_o ? n4890_o : n5333_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5411_o = n4831_o ? n4892_o : n5338_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5412_o = n4831_o ? n4893_o : n5339_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5413_o = n4831_o ? n2148_o : n5340_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5414_o = n4831_o ? n2151_o : n5341_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5415_o = n4831_o ? n4858_o : n5342_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5417_o = n4831_o ? n4896_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5419_o = n4831_o ? n4899_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5421_o = n4831_o ? 1'b0 : n5344_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5423_o = n4831_o ? 1'b0 : n5346_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5424_o = n4831_o ? n1906_o : n5347_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5425_o = n4831_o ? n2154_o : n5348_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5426_o = n4831_o ? n4902_o : n5351_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5428_o = n4831_o ? 1'b0 : n5353_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5430_o = n4831_o ? 1'b0 : n5356_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5432_o = n4831_o ? 1'b0 : n5358_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5433_o = n4831_o ? n4905_o : n5362_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5435_o = n4831_o ? 1'b0 : n5364_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5437_o = n4831_o ? n4908_o : 1'b0;
  assign n5438_o = {n5380_o, n5376_o};
  assign n5439_o = {n5388_o, n5386_o};
  assign n5440_o = {n5398_o, n5393_o};
  assign n5441_o = n1909_o[0];
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5442_o = n4831_o ? n5441_o : n5366_o;
  assign n5443_o = n1909_o[24];
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5444_o = n4831_o ? n5443_o : n5368_o;
  assign n5445_o = n1909_o[34];
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5446_o = n4831_o ? n5445_o : n5370_o;
  assign n5447_o = n1909_o[44];
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5448_o = n4831_o ? n5447_o : n5372_o;
  assign n5449_o = n5438_o[0];
  assign n5450_o = n2162_o[0];
  assign n5451_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n5452_o = n2037_o ? n5450_o : n5451_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5453_o = n4831_o ? n5452_o : n5449_o;
  assign n5454_o = n5438_o[1];
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5455_o = n4831_o ? n4913_o : n5454_o;
  assign n5456_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5457_o = n4831_o ? n5456_o : n5382_o;
  assign n5458_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5459_o = n4831_o ? n5458_o : n5384_o;
  assign n5460_o = n1909_o[60:57];
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5461_o = n4831_o ? n5460_o : n5439_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5462_o = n4844_o & n4831_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5463_o = n4831_o ? n2019_o : n5440_o;
  assign n5464_o = n1909_o[74];
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5465_o = n4831_o ? n5464_o : n5400_o;
  assign n5466_o = {n5408_o, n5406_o};
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5468_o = n4831_o ? 1'b0 : n5402_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5470_o = n4831_o ? 1'b0 : n5404_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5472_o = n4831_o ? 3'b000 : n5466_o;
  /* TG68KdotC_Kernel.vhd:2433:57  */
  assign n5473_o = n4831_o ? n4915_o : n5409_o;
  /* TG68KdotC_Kernel.vhd:2415:49  */
  assign n5475_o = n3613_o == 3'b111;
  assign n5476_o = {n5475_o, n4830_o, n4720_o, n4016_o, n3876_o, n3769_o, n3700_o};
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5477_o = n5410_o;
      7'b0100000: n5477_o = make_berr;
      7'b0010000: n5477_o = make_berr;
      7'b0001000: n5477_o = make_berr;
      7'b0000100: n5477_o = make_berr;
      7'b0000010: n5477_o = n3753_o;
      7'b0000001: n5477_o = n3636_o;
      default: n5477_o = make_berr;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5478_o = n5411_o;
      7'b0100000: n5478_o = n4810_o;
      7'b0010000: n5478_o = n4643_o;
      7'b0001000: n5478_o = n3921_o;
      7'b0000100: n5478_o = n3798_o;
      7'b0000010: n5478_o = n1921_o;
      7'b0000001: n5478_o = n3657_o;
      default: n5478_o = n1921_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5479_o = n5412_o;
      7'b0100000: n5479_o = n2026_o;
      7'b0010000: n5479_o = n4644_o;
      7'b0001000: n5479_o = n3919_o;
      7'b0000100: n5479_o = n2026_o;
      7'b0000010: n5479_o = n2026_o;
      7'b0000001: n5479_o = n2026_o;
      default: n5479_o = n2026_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5480_o = n5413_o;
      7'b0100000: n5480_o = n2148_o;
      7'b0010000: n5480_o = n2148_o;
      7'b0001000: n5480_o = n2148_o;
      7'b0000100: n5480_o = n2148_o;
      7'b0000010: n5480_o = n2148_o;
      7'b0000001: n5480_o = n2148_o;
      default: n5480_o = n2148_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5481_o = n5414_o;
      7'b0100000: n5481_o = n2151_o;
      7'b0010000: n5481_o = n2151_o;
      7'b0001000: n5481_o = n2151_o;
      7'b0000100: n5481_o = n2151_o;
      7'b0000010: n5481_o = n2151_o;
      7'b0000001: n5481_o = n2151_o;
      default: n5481_o = n2151_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5483_o = 1'b0;
      7'b0100000: n5483_o = n4812_o;
      7'b0010000: n5483_o = n4646_o;
      7'b0001000: n5483_o = n3997_o;
      7'b0000100: n5483_o = n3860_o;
      7'b0000010: n5483_o = n3755_o;
      7'b0000001: n5483_o = n3676_o;
      default: n5483_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5484_o = n5415_o;
      7'b0100000: n5484_o = n2015_o;
      7'b0010000: n5484_o = n4647_o;
      7'b0001000: n5484_o = n2015_o;
      7'b0000100: n5484_o = n2015_o;
      7'b0000010: n5484_o = n2015_o;
      7'b0000001: n5484_o = n2015_o;
      default: n5484_o = n2015_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5486_o = n5417_o;
      7'b0100000: n5486_o = 1'b0;
      7'b0010000: n5486_o = 1'b0;
      7'b0001000: n5486_o = 1'b0;
      7'b0000100: n5486_o = 1'b0;
      7'b0000010: n5486_o = 1'b0;
      7'b0000001: n5486_o = 1'b0;
      default: n5486_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5488_o = 1'b0;
      7'b0100000: n5488_o = n4814_o;
      7'b0010000: n5488_o = 1'b0;
      7'b0001000: n5488_o = 1'b0;
      7'b0000100: n5488_o = 1'b0;
      7'b0000010: n5488_o = 1'b0;
      7'b0000001: n5488_o = 1'b0;
      default: n5488_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5490_o = n5419_o;
      7'b0100000: n5490_o = 1'b0;
      7'b0010000: n5490_o = n4648_o;
      7'b0001000: n5490_o = 1'b0;
      7'b0000100: n5490_o = 1'b0;
      7'b0000010: n5490_o = 1'b0;
      7'b0000001: n5490_o = 1'b0;
      default: n5490_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5492_o = n5421_o;
      7'b0100000: n5492_o = n4816_o;
      7'b0010000: n5492_o = n4650_o;
      7'b0001000: n5492_o = 1'b0;
      7'b0000100: n5492_o = 1'b0;
      7'b0000010: n5492_o = 1'b0;
      7'b0000001: n5492_o = 1'b0;
      default: n5492_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5494_o = n5423_o;
      7'b0100000: n5494_o = n4818_o;
      7'b0010000: n5494_o = n4651_o;
      7'b0001000: n5494_o = n3999_o;
      7'b0000100: n5494_o = n3861_o;
      7'b0000010: n5494_o = 1'b0;
      7'b0000001: n5494_o = n3678_o;
      default: n5494_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5496_o = 1'b0;
      7'b0100000: n5496_o = 1'b0;
      7'b0010000: n5496_o = n4653_o;
      7'b0001000: n5496_o = 1'b0;
      7'b0000100: n5496_o = 1'b0;
      7'b0000010: n5496_o = 1'b0;
      7'b0000001: n5496_o = 1'b0;
      default: n5496_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5498_o = 1'b0;
      7'b0100000: n5498_o = 1'b0;
      7'b0010000: n5498_o = n4655_o;
      7'b0001000: n5498_o = 1'b0;
      7'b0000100: n5498_o = 1'b0;
      7'b0000010: n5498_o = 1'b0;
      7'b0000001: n5498_o = 1'b0;
      default: n5498_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5500_o = 1'b0;
      7'b0100000: n5500_o = 1'b0;
      7'b0010000: n5500_o = n4657_o;
      7'b0001000: n5500_o = 1'b0;
      7'b0000100: n5500_o = 1'b0;
      7'b0000010: n5500_o = 1'b0;
      7'b0000001: n5500_o = 1'b0;
      default: n5500_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5501_o = n5424_o;
      7'b0100000: n5501_o = n1906_o;
      7'b0010000: n5501_o = n1906_o;
      7'b0001000: n5501_o = n1906_o;
      7'b0000100: n5501_o = n1906_o;
      7'b0000010: n5501_o = n1906_o;
      7'b0000001: n5501_o = n1906_o;
      default: n5501_o = n1906_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5503_o = 1'b0;
      7'b0100000: n5503_o = 1'b0;
      7'b0010000: n5503_o = n4659_o;
      7'b0001000: n5503_o = 1'b0;
      7'b0000100: n5503_o = 1'b0;
      7'b0000010: n5503_o = 1'b0;
      7'b0000001: n5503_o = 1'b0;
      default: n5503_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5504_o = n5425_o;
      7'b0100000: n5504_o = n2154_o;
      7'b0010000: n5504_o = n2154_o;
      7'b0001000: n5504_o = n2154_o;
      7'b0000100: n5504_o = n2154_o;
      7'b0000010: n5504_o = n2154_o;
      7'b0000001: n5504_o = n2154_o;
      default: n5504_o = n2154_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5506_o = n5426_o;
      7'b0100000: n5506_o = n4820_o;
      7'b0010000: n5506_o = n4660_o;
      7'b0001000: n5506_o = n4000_o;
      7'b0000100: n5506_o = n3862_o;
      7'b0000010: n5506_o = n3757_o;
      7'b0000001: n5506_o = n3681_o;
      default: n5506_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5508_o = n5428_o;
      7'b0100000: n5508_o = 1'b0;
      7'b0010000: n5508_o = 1'b0;
      7'b0001000: n5508_o = n4002_o;
      7'b0000100: n5508_o = 1'b0;
      7'b0000010: n5508_o = 1'b0;
      7'b0000001: n5508_o = 1'b0;
      default: n5508_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5510_o = n5430_o;
      7'b0100000: n5510_o = 1'b0;
      7'b0010000: n5510_o = 1'b0;
      7'b0001000: n5510_o = 1'b0;
      7'b0000100: n5510_o = 1'b0;
      7'b0000010: n5510_o = 1'b0;
      7'b0000001: n5510_o = 1'b0;
      default: n5510_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5512_o = n5432_o;
      7'b0100000: n5512_o = 1'b0;
      7'b0010000: n5512_o = 1'b0;
      7'b0001000: n5512_o = 1'b0;
      7'b0000100: n5512_o = 1'b0;
      7'b0000010: n5512_o = 1'b0;
      7'b0000001: n5512_o = 1'b0;
      default: n5512_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5514_o = n5433_o;
      7'b0100000: n5514_o = n4822_o;
      7'b0010000: n5514_o = n4661_o;
      7'b0001000: n5514_o = n4003_o;
      7'b0000100: n5514_o = n3863_o;
      7'b0000010: n5514_o = n3759_o;
      7'b0000001: n5514_o = n3684_o;
      default: n5514_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5516_o = n5435_o;
      7'b0100000: n5516_o = 1'b0;
      7'b0010000: n5516_o = 1'b0;
      7'b0001000: n5516_o = 1'b0;
      7'b0000100: n5516_o = 1'b0;
      7'b0000010: n5516_o = 1'b0;
      7'b0000001: n5516_o = 1'b0;
      default: n5516_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5518_o = n5437_o;
      7'b0100000: n5518_o = n4824_o;
      7'b0010000: n5518_o = n4663_o;
      7'b0001000: n5518_o = n4004_o;
      7'b0000100: n5518_o = n3864_o;
      7'b0000010: n5518_o = n3761_o;
      7'b0000001: n5518_o = n3687_o;
      default: n5518_o = 1'b0;
    endcase
  assign n5519_o = n1909_o[0];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5520_o = n5442_o;
      7'b0100000: n5520_o = n5519_o;
      7'b0010000: n5520_o = n4665_o;
      7'b0001000: n5520_o = n5519_o;
      7'b0000100: n5520_o = n5519_o;
      7'b0000010: n5520_o = n5519_o;
      7'b0000001: n5520_o = n5519_o;
      default: n5520_o = n5519_o;
    endcase
  assign n5521_o = n1909_o[24];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5522_o = n5444_o;
      7'b0100000: n5522_o = n5521_o;
      7'b0010000: n5522_o = n4667_o;
      7'b0001000: n5522_o = n5521_o;
      7'b0000100: n5522_o = n5521_o;
      7'b0000010: n5522_o = n5521_o;
      7'b0000001: n5522_o = n5521_o;
      default: n5522_o = n5521_o;
    endcase
  assign n5523_o = n1909_o[34];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5524_o = n5446_o;
      7'b0100000: n5524_o = n5523_o;
      7'b0010000: n5524_o = n4669_o;
      7'b0001000: n5524_o = n5523_o;
      7'b0000100: n5524_o = n5523_o;
      7'b0000010: n5524_o = n5523_o;
      7'b0000001: n5524_o = n5523_o;
      default: n5524_o = n5523_o;
    endcase
  assign n5525_o = n1909_o[36];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5526_o = n5525_o;
      7'b0100000: n5526_o = n5525_o;
      7'b0010000: n5526_o = n4671_o;
      7'b0001000: n5526_o = n5525_o;
      7'b0000100: n5526_o = n5525_o;
      7'b0000010: n5526_o = n5525_o;
      7'b0000001: n5526_o = n5525_o;
      default: n5526_o = n5525_o;
    endcase
  assign n5527_o = n1909_o[40];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5528_o = n5527_o;
      7'b0100000: n5528_o = n5527_o;
      7'b0010000: n5528_o = n4673_o;
      7'b0001000: n5528_o = n5527_o;
      7'b0000100: n5528_o = n5527_o;
      7'b0000010: n5528_o = n5527_o;
      7'b0000001: n5528_o = n5527_o;
      default: n5528_o = n5527_o;
    endcase
  assign n5529_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5530_o = n5529_o;
      7'b0100000: n5530_o = n5529_o;
      7'b0010000: n5530_o = n4674_o;
      7'b0001000: n5530_o = n5529_o;
      7'b0000100: n5530_o = n5529_o;
      7'b0000010: n5530_o = n5529_o;
      7'b0000001: n5530_o = n5529_o;
      default: n5530_o = n5529_o;
    endcase
  assign n5531_o = n1909_o[44];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5532_o = n5448_o;
      7'b0100000: n5532_o = n5531_o;
      7'b0010000: n5532_o = n4676_o;
      7'b0001000: n5532_o = n5531_o;
      7'b0000100: n5532_o = n5531_o;
      7'b0000010: n5532_o = n5531_o;
      7'b0000001: n5532_o = n5531_o;
      default: n5532_o = n5531_o;
    endcase
  assign n5533_o = n2162_o[0];
  assign n5534_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n5535_o = n2037_o ? n5533_o : n5534_o;
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5536_o = n5453_o;
      7'b0100000: n5536_o = n5535_o;
      7'b0010000: n5536_o = n5535_o;
      7'b0001000: n5536_o = n5535_o;
      7'b0000100: n5536_o = n5535_o;
      7'b0000010: n5536_o = n5535_o;
      7'b0000001: n5536_o = n5535_o;
      default: n5536_o = n5535_o;
    endcase
  assign n5537_o = n2162_o[1];
  assign n5538_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n5539_o = n2037_o ? n5537_o : n5538_o;
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5540_o = n5455_o;
      7'b0100000: n5540_o = n5539_o;
      7'b0010000: n5540_o = n4680_o;
      7'b0001000: n5540_o = n5539_o;
      7'b0000100: n5540_o = n5539_o;
      7'b0000010: n5540_o = n5539_o;
      7'b0000001: n5540_o = n5539_o;
      default: n5540_o = n5539_o;
    endcase
  assign n5541_o = n1909_o[48];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5542_o = n5541_o;
      7'b0100000: n5542_o = n5541_o;
      7'b0010000: n5542_o = n4683_o;
      7'b0001000: n5542_o = n5541_o;
      7'b0000100: n5542_o = n5541_o;
      7'b0000010: n5542_o = n5541_o;
      7'b0000001: n5542_o = n5541_o;
      default: n5542_o = n5541_o;
    endcase
  assign n5543_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5544_o = n5457_o;
      7'b0100000: n5544_o = n5543_o;
      7'b0010000: n5544_o = n4685_o;
      7'b0001000: n5544_o = n5543_o;
      7'b0000100: n5544_o = n5543_o;
      7'b0000010: n5544_o = n5543_o;
      7'b0000001: n5544_o = n5543_o;
      default: n5544_o = n5543_o;
    endcase
  assign n5545_o = n3905_o[0];
  assign n5546_o = n1909_o[51];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5547_o = n5546_o;
      7'b0100000: n5547_o = n5546_o;
      7'b0010000: n5547_o = n5546_o;
      7'b0001000: n5547_o = n5545_o;
      7'b0000100: n5547_o = n3796_o;
      7'b0000010: n5547_o = n5546_o;
      7'b0000001: n5547_o = n5546_o;
      default: n5547_o = n5546_o;
    endcase
  assign n5548_o = n3905_o[1];
  assign n5549_o = n1909_o[52];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5550_o = n5549_o;
      7'b0100000: n5550_o = n5549_o;
      7'b0010000: n5550_o = n5549_o;
      7'b0001000: n5550_o = n5548_o;
      7'b0000100: n5550_o = n5549_o;
      7'b0000010: n5550_o = n5549_o;
      7'b0000001: n5550_o = n5549_o;
      default: n5550_o = n5549_o;
    endcase
  assign n5551_o = n1909_o[53];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5552_o = n5551_o;
      7'b0100000: n5552_o = n5551_o;
      7'b0010000: n5552_o = n5551_o;
      7'b0001000: n5552_o = n4008_o;
      7'b0000100: n5552_o = n5551_o;
      7'b0000010: n5552_o = n5551_o;
      7'b0000001: n5552_o = n5551_o;
      default: n5552_o = n5551_o;
    endcase
  assign n5553_o = n1909_o[54];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5554_o = n5553_o;
      7'b0100000: n5554_o = n5553_o;
      7'b0010000: n5554_o = n4688_o;
      7'b0001000: n5554_o = n5553_o;
      7'b0000100: n5554_o = n3868_o;
      7'b0000010: n5554_o = n3763_o;
      7'b0000001: n5554_o = n3689_o;
      default: n5554_o = n5553_o;
    endcase
  assign n5555_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5556_o = n5459_o;
      7'b0100000: n5556_o = n5555_o;
      7'b0010000: n5556_o = n4690_o;
      7'b0001000: n5556_o = n5555_o;
      7'b0000100: n5556_o = n5555_o;
      7'b0000010: n5556_o = n5555_o;
      7'b0000001: n5556_o = n5555_o;
      default: n5556_o = n5555_o;
    endcase
  assign n5557_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5558_o = n5557_o;
      7'b0100000: n5558_o = n5557_o;
      7'b0010000: n5558_o = n4693_o;
      7'b0001000: n5558_o = n5557_o;
      7'b0000100: n5558_o = n3870_o;
      7'b0000010: n5558_o = n5557_o;
      7'b0000001: n5558_o = n3691_o;
      default: n5558_o = n5557_o;
    endcase
  assign n5559_o = n1909_o[60:57];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5560_o = n5461_o;
      7'b0100000: n5560_o = n5559_o;
      7'b0010000: n5560_o = n5559_o;
      7'b0001000: n5560_o = n5559_o;
      7'b0000100: n5560_o = n5559_o;
      7'b0000010: n5560_o = n5559_o;
      7'b0000001: n5560_o = n5559_o;
      default: n5560_o = n5559_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5561_o = n4914_o;
      7'b0100000: n5561_o = n2178_o;
      7'b0010000: n5561_o = n2178_o;
      7'b0001000: n5561_o = n2178_o;
      7'b0000100: n5561_o = n2178_o;
      7'b0000010: n5561_o = n2178_o;
      7'b0000001: n5561_o = n2178_o;
      default: n5561_o = n2178_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5562_o = n5463_o;
      7'b0100000: n5562_o = n2019_o;
      7'b0010000: n5562_o = n2019_o;
      7'b0001000: n5562_o = n2019_o;
      7'b0000100: n5562_o = n2019_o;
      7'b0000010: n5562_o = n2019_o;
      7'b0000001: n5562_o = n2019_o;
      default: n5562_o = n2019_o;
    endcase
  assign n5563_o = n1909_o[69];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5564_o = n5563_o;
      7'b0100000: n5564_o = n5563_o;
      7'b0010000: n5564_o = n4695_o;
      7'b0001000: n5564_o = n5563_o;
      7'b0000100: n5564_o = n5563_o;
      7'b0000010: n5564_o = n5563_o;
      7'b0000001: n5564_o = n5563_o;
      default: n5564_o = n5563_o;
    endcase
  assign n5565_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5566_o = n5565_o;
      7'b0100000: n5566_o = n5565_o;
      7'b0010000: n5566_o = n4696_o;
      7'b0001000: n5566_o = n5565_o;
      7'b0000100: n5566_o = n5565_o;
      7'b0000010: n5566_o = n5565_o;
      7'b0000001: n5566_o = n5565_o;
      default: n5566_o = n5565_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5567_o = n2171_o;
      7'b0100000: n5567_o = n2171_o;
      7'b0010000: n5567_o = n4697_o;
      7'b0001000: n5567_o = n2171_o;
      7'b0000100: n5567_o = n2171_o;
      7'b0000010: n5567_o = n2171_o;
      7'b0000001: n5567_o = n2171_o;
      default: n5567_o = n2171_o;
    endcase
  assign n5568_o = n1909_o[74];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5569_o = n5465_o;
      7'b0100000: n5569_o = n5568_o;
      7'b0010000: n5569_o = n5568_o;
      7'b0001000: n5569_o = n5568_o;
      7'b0000100: n5569_o = n5568_o;
      7'b0000010: n5569_o = n5568_o;
      7'b0000001: n5569_o = n5568_o;
      default: n5569_o = n5568_o;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5571_o = n5468_o;
      7'b0100000: n5571_o = n4826_o;
      7'b0010000: n5571_o = n4699_o;
      7'b0001000: n5571_o = 1'b0;
      7'b0000100: n5571_o = 1'b0;
      7'b0000010: n5571_o = 1'b0;
      7'b0000001: n5571_o = 1'b0;
      default: n5571_o = 1'b0;
    endcase
  assign n5572_o = n3694_o[0];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5574_o = 1'b0;
      7'b0100000: n5574_o = 1'b0;
      7'b0010000: n5574_o = 1'b0;
      7'b0001000: n5574_o = 1'b0;
      7'b0000100: n5574_o = 1'b0;
      7'b0000010: n5574_o = 1'b0;
      7'b0000001: n5574_o = n5572_o;
      default: n5574_o = 1'b0;
    endcase
  assign n5575_o = n3694_o[1];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5577_o = n5470_o;
      7'b0100000: n5577_o = 1'b0;
      7'b0010000: n5577_o = n4701_o;
      7'b0001000: n5577_o = 1'b0;
      7'b0000100: n5577_o = n3872_o;
      7'b0000010: n5577_o = 1'b0;
      7'b0000001: n5577_o = n5575_o;
      default: n5577_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5579_o = 1'b0;
      7'b0100000: n5579_o = 1'b0;
      7'b0010000: n5579_o = 1'b0;
      7'b0001000: n5579_o = 1'b0;
      7'b0000100: n5579_o = 1'b0;
      7'b0000010: n5579_o = n3765_o;
      7'b0000001: n5579_o = 1'b0;
      default: n5579_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5581_o = 1'b0;
      7'b0100000: n5581_o = 1'b0;
      7'b0010000: n5581_o = 1'b0;
      7'b0001000: n5581_o = n4010_o;
      7'b0000100: n5581_o = 1'b0;
      7'b0000010: n5581_o = 1'b0;
      7'b0000001: n5581_o = 1'b0;
      default: n5581_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5583_o = 1'b0;
      7'b0100000: n5583_o = 1'b0;
      7'b0010000: n5583_o = n4703_o;
      7'b0001000: n5583_o = 1'b0;
      7'b0000100: n5583_o = 1'b0;
      7'b0000010: n5583_o = 1'b0;
      7'b0000001: n5583_o = 1'b0;
      default: n5583_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5585_o = 1'b0;
      7'b0100000: n5585_o = 1'b0;
      7'b0010000: n5585_o = n4705_o;
      7'b0001000: n5585_o = 1'b0;
      7'b0000100: n5585_o = 1'b0;
      7'b0000010: n5585_o = 1'b0;
      7'b0000001: n5585_o = 1'b0;
      default: n5585_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5587_o = 1'b0;
      7'b0100000: n5587_o = 1'b0;
      7'b0010000: n5587_o = n4707_o;
      7'b0001000: n5587_o = 1'b0;
      7'b0000100: n5587_o = 1'b0;
      7'b0000010: n5587_o = 1'b0;
      7'b0000001: n5587_o = 1'b0;
      default: n5587_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5589_o = 1'b0;
      7'b0100000: n5589_o = 1'b0;
      7'b0010000: n5589_o = 1'b0;
      7'b0001000: n5589_o = n4012_o;
      7'b0000100: n5589_o = 1'b0;
      7'b0000010: n5589_o = 1'b0;
      7'b0000001: n5589_o = 1'b0;
      default: n5589_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5591_o = 1'b0;
      7'b0100000: n5591_o = 1'b0;
      7'b0010000: n5591_o = n4709_o;
      7'b0001000: n5591_o = 1'b0;
      7'b0000100: n5591_o = 1'b0;
      7'b0000010: n5591_o = 1'b0;
      7'b0000001: n5591_o = n3696_o;
      default: n5591_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5593_o = 1'b0;
      7'b0100000: n5593_o = 1'b0;
      7'b0010000: n5593_o = n4711_o;
      7'b0001000: n5593_o = 1'b0;
      7'b0000100: n5593_o = 1'b0;
      7'b0000010: n5593_o = 1'b0;
      7'b0000001: n5593_o = 1'b0;
      default: n5593_o = 1'b0;
    endcase
  assign n5594_o = n5472_o[1:0];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5596_o = n5594_o;
      7'b0100000: n5596_o = 2'b00;
      7'b0010000: n5596_o = 2'b00;
      7'b0001000: n5596_o = 2'b00;
      7'b0000100: n5596_o = 2'b00;
      7'b0000010: n5596_o = 2'b00;
      7'b0000001: n5596_o = 2'b00;
      default: n5596_o = 2'b00;
    endcase
  assign n5597_o = n5472_o[2];
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5599_o = n5597_o;
      7'b0100000: n5599_o = n4828_o;
      7'b0010000: n5599_o = n4712_o;
      7'b0001000: n5599_o = n4014_o;
      7'b0000100: n5599_o = n3874_o;
      7'b0000010: n5599_o = n3767_o;
      7'b0000001: n5599_o = n3698_o;
      default: n5599_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5601_o = 1'b0;
      7'b0100000: n5601_o = 1'b0;
      7'b0010000: n5601_o = n4714_o;
      7'b0001000: n5601_o = 1'b0;
      7'b0000100: n5601_o = 1'b0;
      7'b0000010: n5601_o = 1'b0;
      7'b0000001: n5601_o = 1'b0;
      default: n5601_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:2044:41  */
  always @*
    case (n5476_o)
      7'b1000000: n5602_o = n5473_o;
      7'b0100000: n5602_o = n2180_o;
      7'b0010000: n5602_o = n4715_o;
      7'b0001000: n5602_o = n2180_o;
      7'b0000100: n5602_o = n2180_o;
      7'b0000010: n5602_o = n2180_o;
      7'b0000001: n5602_o = n2180_o;
      default: n5602_o = n2180_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5603_o = n3356_o ? make_berr : n5477_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5604_o = n3356_o ? n3583_o : n5478_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5605_o = n3356_o ? n3584_o : n5479_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5606_o = n3356_o ? n2148_o : n5480_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5607_o = n3356_o ? n2151_o : n5481_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5609_o = n3356_o ? 1'b0 : n5483_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5610_o = n3356_o ? n2015_o : n5484_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5612_o = n3356_o ? 1'b0 : n5486_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5614_o = n3356_o ? 1'b0 : n5488_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5615_o = n3356_o ? n3586_o : n5490_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5616_o = n3356_o ? n3588_o : n5492_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5617_o = n3356_o ? n3589_o : n5494_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5619_o = n3356_o ? 1'b0 : n5496_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5621_o = n3356_o ? n3591_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5623_o = n3356_o ? 1'b0 : n5498_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5624_o = n3356_o ? n3592_o : n5500_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5625_o = n3356_o ? n1906_o : n5501_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5627_o = n3356_o ? 1'b0 : n5503_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5628_o = n3356_o ? n3593_o : n5504_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5629_o = n3356_o ? n3594_o : n5506_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5631_o = n3356_o ? 1'b0 : n5508_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5633_o = n3356_o ? 1'b0 : n5510_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5635_o = n3356_o ? 1'b0 : n5512_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5636_o = n3356_o ? n3595_o : n5514_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5638_o = n3356_o ? 1'b0 : n5516_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5639_o = n3356_o ? n3596_o : n5518_o;
  assign n5640_o = {n5544_o, n5542_o, n5540_o, n5536_o};
  assign n5641_o = {n5560_o, n5558_o, n5556_o, n5554_o, n5552_o, n5550_o, n5547_o};
  assign n5642_o = {n5562_o, n5561_o};
  assign n5643_o = {n5569_o, n5567_o};
  assign n5644_o = n1909_o[0];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5645_o = n3356_o ? n5644_o : n5520_o;
  assign n5646_o = n1909_o[24];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5647_o = n3356_o ? n5646_o : n5522_o;
  assign n5648_o = n1909_o[34];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5649_o = n3356_o ? n5648_o : n5524_o;
  assign n5650_o = n1909_o[36];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5651_o = n3356_o ? n5650_o : n5526_o;
  assign n5652_o = n1909_o[40];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5653_o = n3356_o ? n5652_o : n5528_o;
  assign n5654_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5655_o = n3356_o ? n5654_o : n5530_o;
  assign n5656_o = n1909_o[43];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5657_o = n3356_o ? n3598_o : n5656_o;
  assign n5658_o = n1909_o[44];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5659_o = n3356_o ? n5658_o : n5532_o;
  assign n5660_o = n5640_o[2:0];
  assign n5661_o = n1909_o[48];
  assign n5662_o = {n5661_o, n2166_o};
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5663_o = n3356_o ? n5662_o : n5660_o;
  assign n5664_o = n5640_o[3];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5665_o = n3356_o ? n3600_o : n5664_o;
  assign n5666_o = n5641_o[4:0];
  assign n5667_o = n1909_o[55:51];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5668_o = n3356_o ? n5667_o : n5666_o;
  assign n5669_o = n5641_o[5];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5670_o = n3356_o ? n3602_o : n5669_o;
  assign n5671_o = n5641_o[9:6];
  assign n5672_o = n1909_o[60:57];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5673_o = n3356_o ? n5672_o : n5671_o;
  assign n5674_o = {n2019_o, n2178_o};
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5675_o = n3356_o ? n5674_o : n5642_o;
  assign n5676_o = n1909_o[69];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5677_o = n3356_o ? n5676_o : n5564_o;
  assign n5678_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5679_o = n3356_o ? n5678_o : n5566_o;
  assign n5680_o = n1909_o[74];
  assign n5681_o = {n5680_o, n2171_o};
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5682_o = n3356_o ? n5681_o : n5643_o;
  assign n5683_o = {n5577_o, n5574_o};
  assign n5684_o = {n5581_o, n5579_o};
  assign n5685_o = {n5599_o, n5596_o};
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5686_o = n3356_o ? n3604_o : n5571_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5688_o = n3356_o ? 2'b00 : n5683_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5690_o = n3356_o ? 2'b00 : n5684_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5691_o = n3356_o ? n3606_o : n5583_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5693_o = n3356_o ? 1'b0 : n5585_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5695_o = n3356_o ? 1'b0 : n5587_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5697_o = n3356_o ? 1'b0 : n5589_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5699_o = n3356_o ? 1'b0 : n5591_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5701_o = n3356_o ? 1'b0 : n5593_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5703_o = n3356_o ? n3608_o : 1'b0;
  assign n5704_o = n5685_o[1:0];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5706_o = n3356_o ? 2'b00 : n5704_o;
  assign n5707_o = n5685_o[2];
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5708_o = n3356_o ? n3610_o : n5707_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5709_o = n3356_o ? n3612_o : n5601_o;
  /* TG68KdotC_Kernel.vhd:1966:33  */
  assign n5710_o = n3356_o ? n2180_o : n5602_o;
  /* TG68KdotC_Kernel.vhd:1965:25  */
  assign n5712_o = n2185_o == 4'b0100;
  /* TG68KdotC_Kernel.vhd:2644:50  */
  assign n5713_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2644:62  */
  assign n5715_o = n5713_o == 2'b11;
  /* TG68KdotC_Kernel.vhd:2645:58  */
  assign n5716_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2645:70  */
  assign n5718_o = n5716_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:2646:57  */
  assign n5722_o = decodeopc ? 1'b1 : 1'b0;
  assign n5723_o = n1909_o[53];
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n5724_o = n5919_o ? 1'b1 : n5723_o;
  /* TG68KdotC_Kernel.vhd:2646:57  */
  assign n5726_o = decodeopc ? 7'b0011001 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2651:61  */
  assign n5727_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2651:73  */
  assign n5729_o = n5727_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:2651:91  */
  assign n5730_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2651:103  */
  assign n5732_o = n5730_o == 2'b01;
  /* TG68KdotC_Kernel.vhd:2651:118  */
  assign n5733_o = opcode[2:0];
  /* TG68KdotC_Kernel.vhd:2651:130  */
  assign n5735_o = n5733_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:2651:109  */
  assign n5736_o = n5732_o | n5735_o;
  /* TG68KdotC_Kernel.vhd:2651:80  */
  assign n5737_o = n5736_o & n5729_o;
  /* TG68KdotC_Kernel.vhd:2652:63  */
  assign n5738_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:2653:74  */
  assign n5739_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2653:86  */
  assign n5741_o = n5739_o == 2'b01;
  /* TG68KdotC_Kernel.vhd:2655:90  */
  assign n5742_o = opcode[0];
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5744_o = n5823_o ? 1'b1 : n2171_o;
  /* TG68KdotC_Kernel.vhd:2654:73  */
  assign n5745_o = n5742_o & decodeopc;
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5747_o = n5828_o ? 7'b0000001 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2661:73  */
  assign n5749_o = decodeopc ? 2'b01 : n2026_o;
  /* TG68KdotC_Kernel.vhd:2653:65  */
  assign n5750_o = n5741_o ? n2026_o : n5749_o;
  /* TG68KdotC_Kernel.vhd:2653:65  */
  assign n5751_o = n5745_o & n5741_o;
  /* TG68KdotC_Kernel.vhd:2653:65  */
  assign n5752_o = decodeopc & n5741_o;
  /* TG68KdotC_Kernel.vhd:2665:99  */
  assign n5753_o = ~decodeopc;
  /* TG68KdotC_Kernel.vhd:2665:86  */
  assign n5754_o = n5753_o & exe_condition;
  /* TG68KdotC_Kernel.vhd:2665:65  */
  assign n5757_o = n5754_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2665:65  */
  assign n5760_o = n5754_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5761_o = n5814_o ? n5750_o : n2026_o;
  /* TG68KdotC_Kernel.vhd:2652:57  */
  assign n5764_o = n5738_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2652:57  */
  assign n5766_o = n5738_o ? n5757_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2652:57  */
  assign n5768_o = n5738_o ? n5760_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:2652:57  */
  assign n5769_o = n5751_o & n5738_o;
  /* TG68KdotC_Kernel.vhd:2652:57  */
  assign n5770_o = n5752_o & n5738_o;
  /* TG68KdotC_Kernel.vhd:2673:62  */
  assign n5771_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2673:74  */
  assign n5773_o = n5771_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:2673:91  */
  assign n5774_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2673:103  */
  assign n5776_o = n5774_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2673:82  */
  assign n5777_o = n5773_o | n5776_o;
  /* TG68KdotC_Kernel.vhd:2678:63  */
  assign n5779_o = cpu[0];
  /* TG68KdotC_Kernel.vhd:2678:80  */
  assign n5781_o = state == 2'b10;
  /* TG68KdotC_Kernel.vhd:2678:71  */
  assign n5782_o = n5781_o & n5779_o;
  /* TG68KdotC_Kernel.vhd:2678:99  */
  assign n5783_o = ~addrvalue;
  /* TG68KdotC_Kernel.vhd:2678:86  */
  assign n5784_o = n5783_o & n5782_o;
  /* TG68KdotC_Kernel.vhd:2673:49  */
  assign n5786_o = n5793_o ? 1'b1 : make_berr;
  /* TG68KdotC_Kernel.vhd:2681:66  */
  assign n5787_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2681:78  */
  assign n5789_o = n5787_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2681:57  */
  assign n5792_o = n5789_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2673:49  */
  assign n5793_o = n5784_o & n5777_o;
  /* TG68KdotC_Kernel.vhd:2673:49  */
  assign n5795_o = n5777_o ? 2'b00 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2673:49  */
  assign n5798_o = n5777_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2673:49  */
  assign n5801_o = n5777_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2673:49  */
  assign n5804_o = n5777_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2673:49  */
  assign n5807_o = n5777_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2673:49  */
  assign n5809_o = n5777_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2673:49  */
  assign n5811_o = n5777_o ? n5792_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5812_o = n5737_o ? make_berr : n5786_o;
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5813_o = n5737_o ? n1921_o : n5795_o;
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5814_o = n5738_o & n5737_o;
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5816_o = n5737_o ? 1'b0 : n5798_o;
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5817_o = n5737_o ? n5764_o : n5801_o;
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5819_o = n5737_o ? n5766_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5820_o = n5737_o ? n5768_o : n5804_o;
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5822_o = n5737_o ? 1'b0 : n5807_o;
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5823_o = n5769_o & n5737_o;
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5825_o = n5737_o ? 1'b0 : n5809_o;
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5827_o = n5737_o ? 1'b0 : n5811_o;
  /* TG68KdotC_Kernel.vhd:2651:49  */
  assign n5828_o = n5770_o & n5737_o;
  /* TG68KdotC_Kernel.vhd:2645:49  */
  assign n5829_o = n5718_o ? make_berr : n5812_o;
  /* TG68KdotC_Kernel.vhd:2645:49  */
  assign n5830_o = n5718_o ? n1921_o : n5813_o;
  /* TG68KdotC_Kernel.vhd:2645:49  */
  assign n5831_o = n5718_o ? n2026_o : n5761_o;
  /* TG68KdotC_Kernel.vhd:2645:49  */
  assign n5833_o = n5718_o ? n5722_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2645:49  */
  assign n5835_o = n5718_o ? 1'b0 : n5816_o;
  /* TG68KdotC_Kernel.vhd:2645:49  */
  assign n5837_o = n5718_o ? 1'b0 : n5817_o;
  /* TG68KdotC_Kernel.vhd:2645:49  */
  assign n5839_o = n5718_o ? 1'b0 : n5819_o;
  /* TG68KdotC_Kernel.vhd:2645:49  */
  assign n5841_o = n5718_o ? 1'b0 : n5820_o;
  /* TG68KdotC_Kernel.vhd:2645:49  */
  assign n5843_o = n5718_o ? 1'b0 : n5822_o;
  /* TG68KdotC_Kernel.vhd:2645:49  */
  assign n5845_o = decodeopc & n5718_o;
  /* TG68KdotC_Kernel.vhd:2645:49  */
  assign n5846_o = n5718_o ? n2171_o : n5744_o;
  /* TG68KdotC_Kernel.vhd:2645:49  */
  assign n5848_o = n5718_o ? 1'b0 : n5825_o;
  /* TG68KdotC_Kernel.vhd:2645:49  */
  assign n5850_o = n5718_o ? 1'b0 : n5827_o;
  /* TG68KdotC_Kernel.vhd:2645:49  */
  assign n5851_o = n5718_o ? n5726_o : n5747_o;
  /* TG68KdotC_Kernel.vhd:2689:58  */
  assign n5852_o = opcode[7:3];
  /* TG68KdotC_Kernel.vhd:2689:70  */
  assign n5854_o = n5852_o != 5'b00001;
  /* TG68KdotC_Kernel.vhd:2690:59  */
  assign n5855_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2690:71  */
  assign n5857_o = n5855_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:2690:88  */
  assign n5858_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2690:100  */
  assign n5860_o = n5858_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2690:79  */
  assign n5861_o = n5857_o | n5860_o;
  /* TG68KdotC_Kernel.vhd:2689:80  */
  assign n5862_o = n5861_o & n5854_o;
  /* TG68KdotC_Kernel.vhd:2692:66  */
  assign n5863_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2692:78  */
  assign n5865_o = n5863_o == 3'b001;
  assign n5867_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:2689:49  */
  assign n5868_o = n5895_o ? 1'b1 : n5867_o;
  /* TG68KdotC_Kernel.vhd:2695:66  */
  assign n5869_o = opcode[8];
  assign n5871_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2689:49  */
  assign n5872_o = n5897_o ? 1'b1 : n5871_o;
  /* TG68KdotC_Kernel.vhd:2702:66  */
  assign n5876_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2702:78  */
  assign n5878_o = n5876_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2702:57  */
  assign n5881_o = n5878_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2689:49  */
  assign n5884_o = n5862_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2689:49  */
  assign n5887_o = n5862_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2689:49  */
  assign n5890_o = n5862_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2689:49  */
  assign n5893_o = n5862_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2689:49  */
  assign n5895_o = n5865_o & n5862_o;
  /* TG68KdotC_Kernel.vhd:2689:49  */
  assign n5897_o = n5869_o & n5862_o;
  assign n5898_o = {1'b1, 1'b1};
  /* TG68KdotC_Kernel.vhd:2689:49  */
  assign n5900_o = n5862_o ? n5898_o : 2'b00;
  /* TG68KdotC_Kernel.vhd:2689:49  */
  assign n5902_o = n5862_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2689:49  */
  assign n5904_o = n5862_o ? n5881_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n5905_o = n5715_o ? n5829_o : make_berr;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n5906_o = n5715_o ? n5830_o : n1921_o;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n5907_o = n5715_o ? n5831_o : n2026_o;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n5909_o = n5715_o ? n5833_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n5910_o = n5715_o ? n5835_o : n5884_o;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n5911_o = n5715_o ? n5837_o : n5887_o;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n5913_o = n5715_o ? n5839_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n5914_o = n5715_o ? n5841_o : n5890_o;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n5915_o = n5715_o ? n5843_o : n5893_o;
  assign n5916_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n5917_o = n5715_o ? n5916_o : n5868_o;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n5919_o = n5845_o & n5715_o;
  assign n5920_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n5921_o = n5715_o ? n5920_o : n5872_o;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n5922_o = n5715_o ? n5846_o : n2171_o;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n5924_o = n5715_o ? 2'b00 : n5900_o;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n5926_o = n5715_o ? n5848_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n5928_o = n5715_o ? 1'b0 : n5902_o;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n5929_o = n5715_o ? n5850_o : n5904_o;
  /* TG68KdotC_Kernel.vhd:2644:41  */
  assign n5930_o = n5715_o ? n5851_o : n2180_o;
  /* TG68KdotC_Kernel.vhd:2643:25  */
  assign n5932_o = n2185_o == 4'b0101;
  /* TG68KdotC_Kernel.vhd:2715:47  */
  assign n5934_o = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:2716:50  */
  assign n5935_o = opcode[11:8];
  /* TG68KdotC_Kernel.vhd:2716:63  */
  assign n5937_o = n5935_o == 4'b0001;
  /* TG68KdotC_Kernel.vhd:2719:58  */
  assign n5939_o = opcode[7:0];
  /* TG68KdotC_Kernel.vhd:2719:70  */
  assign n5941_o = n5939_o == 8'b11111111;
  /* TG68KdotC_Kernel.vhd:2722:61  */
  assign n5943_o = opcode[7:0];
  /* TG68KdotC_Kernel.vhd:2722:73  */
  assign n5945_o = n5943_o == 8'b00000000;
  /* TG68KdotC_Kernel.vhd:2722:49  */
  assign n5947_o = n5945_o ? n2026_o : 2'b11;
  /* TG68KdotC_Kernel.vhd:2722:49  */
  assign n5950_o = n5945_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2722:49  */
  assign n5953_o = n5945_o ? 7'b0010111 : 7'b0010110;
  /* TG68KdotC_Kernel.vhd:2719:49  */
  assign n5954_o = n5941_o ? n2026_o : n5947_o;
  /* TG68KdotC_Kernel.vhd:2719:49  */
  assign n5956_o = n5941_o ? 1'b0 : n5950_o;
  /* TG68KdotC_Kernel.vhd:2719:49  */
  assign n5957_o = n5941_o ? 1'b1 : n2171_o;
  /* TG68KdotC_Kernel.vhd:2719:49  */
  assign n5959_o = n5941_o ? 7'b0010111 : n5953_o;
  /* TG68KdotC_Kernel.vhd:2730:58  */
  assign n5960_o = opcode[7:0];
  /* TG68KdotC_Kernel.vhd:2730:70  */
  assign n5962_o = n5960_o == 8'b11111111;
  /* TG68KdotC_Kernel.vhd:2733:61  */
  assign n5964_o = opcode[7:0];
  /* TG68KdotC_Kernel.vhd:2733:73  */
  assign n5966_o = n5964_o == 8'b00000000;
  /* TG68KdotC_Kernel.vhd:2733:49  */
  assign n5968_o = n5966_o ? n2026_o : 2'b01;
  /* TG68KdotC_Kernel.vhd:2730:49  */
  assign n5969_o = n5962_o ? n2026_o : n5968_o;
  /* TG68KdotC_Kernel.vhd:2730:49  */
  assign n5970_o = n5962_o ? 1'b1 : n2171_o;
  /* TG68KdotC_Kernel.vhd:2716:41  */
  assign n5971_o = n5937_o ? n5954_o : n5969_o;
  /* TG68KdotC_Kernel.vhd:2715:33  */
  assign n5973_o = n5984_o ? 1'b1 : n2015_o;
  /* TG68KdotC_Kernel.vhd:2716:41  */
  assign n5975_o = n5937_o ? n5956_o : 1'b0;
  assign n5976_o = n2162_o[1];
  assign n5977_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n5978_o = n2037_o ? n5976_o : n5977_o;
  /* TG68KdotC_Kernel.vhd:2716:41  */
  assign n5979_o = n5937_o ? 1'b1 : n5978_o;
  /* TG68KdotC_Kernel.vhd:2716:41  */
  assign n5980_o = n5937_o ? n5957_o : n5970_o;
  /* TG68KdotC_Kernel.vhd:2716:41  */
  assign n5982_o = n5937_o ? n5959_o : 7'b0010101;
  /* TG68KdotC_Kernel.vhd:2715:33  */
  assign n5983_o = n5934_o ? n5971_o : n2026_o;
  /* TG68KdotC_Kernel.vhd:2715:33  */
  assign n5984_o = n5937_o & n5934_o;
  /* TG68KdotC_Kernel.vhd:2715:33  */
  assign n5986_o = n5934_o ? n5975_o : 1'b0;
  assign n5987_o = n2162_o[1];
  assign n5988_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n5989_o = n2037_o ? n5987_o : n5988_o;
  /* TG68KdotC_Kernel.vhd:2715:33  */
  assign n5990_o = n5934_o ? n5979_o : n5989_o;
  /* TG68KdotC_Kernel.vhd:2715:33  */
  assign n5991_o = n5934_o ? n5980_o : n2171_o;
  /* TG68KdotC_Kernel.vhd:2715:33  */
  assign n5992_o = n5934_o ? n5982_o : n2180_o;
  /* TG68KdotC_Kernel.vhd:2712:25  */
  assign n5994_o = n2185_o == 4'b0110;
  /* TG68KdotC_Kernel.vhd:2744:42  */
  assign n5995_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:2744:45  */
  assign n5996_o = ~n5995_o;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6001_o = n5996_o ? 2'b10 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6004_o = n5996_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6007_o = n5996_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6010_o = n5996_o ? 1'b0 : 1'b1;
  assign n6011_o = {1'b1, 1'b1};
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6013_o = n5996_o ? n6011_o : 2'b00;
  /* TG68KdotC_Kernel.vhd:2744:33  */
  assign n6015_o = n5996_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2743:25  */
  assign n6017_o = n2185_o == 4'b0111;
  /* TG68KdotC_Kernel.vhd:2757:42  */
  assign n6018_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2757:54  */
  assign n6020_o = n6018_o == 2'b11;
  /* TG68KdotC_Kernel.vhd:2759:50  */
  assign n6021_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2759:62  */
  assign n6023_o = n6021_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2758:56  */
  assign n6025_o = n6023_o & 1'b1;
  /* TG68KdotC_Kernel.vhd:2759:81  */
  assign n6026_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2759:93  */
  assign n6028_o = n6026_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2759:111  */
  assign n6029_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:2759:123  */
  assign n6031_o = n6029_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2759:102  */
  assign n6032_o = n6028_o | n6031_o;
  /* TG68KdotC_Kernel.vhd:2759:70  */
  assign n6033_o = n6032_o & n6025_o;
  /* TG68KdotC_Kernel.vhd:2760:58  */
  assign n6034_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2760:70  */
  assign n6036_o = n6034_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2760:49  */
  assign n6039_o = n6036_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2763:64  */
  assign n6041_o = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:2763:70  */
  assign n6042_o = nextpass & n6041_o;
  /* TG68KdotC_Kernel.vhd:2763:98  */
  assign n6043_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2763:110  */
  assign n6045_o = n6043_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2763:116  */
  assign n6046_o = decodeopc & n6045_o;
  /* TG68KdotC_Kernel.vhd:2763:88  */
  assign n6047_o = n6042_o | n6046_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6049_o = n6303_o ? 2'b01 : n2026_o;
  /* TG68KdotC_Kernel.vhd:2758:41  */
  assign n6051_o = n6087_o ? 7'b1011001 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2768:59  */
  assign n6052_o = ~z_error;
  /* TG68KdotC_Kernel.vhd:2768:78  */
  assign n6053_o = ~set_v_flag;
  /* TG68KdotC_Kernel.vhd:2768:64  */
  assign n6054_o = n6053_o & n6052_o;
  /* TG68KdotC_Kernel.vhd:2768:49  */
  assign n6057_o = n6054_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2772:75  */
  assign n6058_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2772:87  */
  assign n6060_o = n6058_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2772:93  */
  assign n6061_o = decodeopc & n6060_o;
  /* TG68KdotC_Kernel.vhd:2772:65  */
  assign n6062_o = nextpass | n6061_o;
  /* TG68KdotC_Kernel.vhd:2772:49  */
  assign n6065_o = n6062_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2758:41  */
  assign n6067_o = n6033_o ? 2'b01 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2758:41  */
  assign n6068_o = n6047_o & n6033_o;
  /* TG68KdotC_Kernel.vhd:2758:41  */
  assign n6070_o = n6033_o ? n6039_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2758:41  */
  assign n6073_o = n6033_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2758:41  */
  assign n6075_o = n6033_o ? n6065_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2758:41  */
  assign n6078_o = n6033_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2758:41  */
  assign n6081_o = n6033_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2758:41  */
  assign n6084_o = n6033_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2758:41  */
  assign n6086_o = n6033_o ? n6057_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2758:41  */
  assign n6087_o = n6047_o & n6033_o;
  /* TG68KdotC_Kernel.vhd:2780:45  */
  assign n6088_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:2780:63  */
  assign n6089_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2780:75  */
  assign n6091_o = n6089_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2780:53  */
  assign n6092_o = n6091_o & n6088_o;
  /* TG68KdotC_Kernel.vhd:2781:50  */
  assign n6093_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2781:62  */
  assign n6095_o = n6093_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2786:53  */
  assign n6099_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2786:65  */
  assign n6101_o = n6099_o == 2'b01;
  /* TG68KdotC_Kernel.vhd:2786:80  */
  assign n6102_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2786:92  */
  assign n6104_o = n6102_o == 2'b10;
  /* TG68KdotC_Kernel.vhd:2786:71  */
  assign n6105_o = n6101_o | n6104_o;
  /* TG68KdotC_Kernel.vhd:2790:58  */
  assign n6108_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2790:71  */
  assign n6110_o = n6108_o == 2'b01;
  /* TG68KdotC_Kernel.vhd:2790:49  */
  assign n6115_o = n6110_o ? 2'b01 : 2'b00;
  /* TG68KdotC_Kernel.vhd:2790:49  */
  assign n6117_o = n6110_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2790:49  */
  assign n6119_o = n6110_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2797:58  */
  assign n6120_o = opcode[3];
  /* TG68KdotC_Kernel.vhd:2797:61  */
  assign n6121_o = ~n6120_o;
  /* TG68KdotC_Kernel.vhd:2798:66  */
  assign n6122_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2798:79  */
  assign n6124_o = n6122_o == 2'b01;
  /* TG68KdotC_Kernel.vhd:2798:57  */
  assign n6127_o = n6124_o ? 2'b00 : 2'b01;
  assign n6131_o = n1909_o[44];
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6132_o = n6173_o ? 1'b1 : n6131_o;
  assign n6133_o = n1909_o[80];
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6134_o = n6177_o ? 1'b1 : n6133_o;
  /* TG68KdotC_Kernel.vhd:2805:57  */
  assign n6136_o = decodeopc ? 7'b0000001 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2813:57  */
  assign n6138_o = decodeopc ? 1'b1 : n2154_o;
  /* TG68KdotC_Kernel.vhd:2813:57  */
  assign n6140_o = decodeopc ? 7'b0011110 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6141_o = n6157_o ? n6127_o : datatype;
  /* TG68KdotC_Kernel.vhd:2797:49  */
  assign n6144_o = n6121_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2797:49  */
  assign n6147_o = n6121_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2797:49  */
  assign n6148_o = n6121_o ? n2154_o : n6138_o;
  /* TG68KdotC_Kernel.vhd:2797:49  */
  assign n6150_o = decodeopc & n6121_o;
  /* TG68KdotC_Kernel.vhd:2797:49  */
  assign n6152_o = decodeopc & n6121_o;
  /* TG68KdotC_Kernel.vhd:2797:49  */
  assign n6154_o = n6121_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2797:49  */
  assign n6155_o = n6121_o ? n6136_o : n6140_o;
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6156_o = n6105_o ? n6115_o : n1921_o;
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6157_o = n6121_o & n6105_o;
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6159_o = n6105_o ? n6144_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6162_o = n6105_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6164_o = n6105_o ? n6147_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6165_o = n6105_o ? n6148_o : n2154_o;
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6168_o = n6105_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6171_o = n6105_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6173_o = n6150_o & n6105_o;
  assign n6174_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6175_o = n6105_o ? 1'b1 : n6174_o;
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6177_o = n6152_o & n6105_o;
  assign n6178_o = {n6119_o, n6117_o};
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6180_o = n6105_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6182_o = n6105_o ? n6154_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6184_o = n6105_o ? n6178_o : 2'b00;
  /* TG68KdotC_Kernel.vhd:2786:41  */
  assign n6185_o = n6105_o ? n6155_o : n2180_o;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6186_o = n6095_o ? n1921_o : n6156_o;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6187_o = n6095_o ? datatype : n6141_o;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6189_o = n6095_o ? 1'b0 : n6159_o;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6191_o = n6095_o ? 1'b0 : n6162_o;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6193_o = n6095_o ? 1'b0 : n6164_o;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6194_o = n6095_o ? n2154_o : n6165_o;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6196_o = n6095_o ? 1'b0 : n6168_o;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6198_o = n6095_o ? 1'b0 : n6171_o;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6201_o = n6095_o ? 1'b1 : 1'b0;
  assign n6202_o = n1909_o[44];
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6203_o = n6095_o ? n6202_o : n6132_o;
  assign n6204_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6205_o = n6095_o ? n6204_o : n6175_o;
  assign n6206_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6207_o = n6285_o ? 1'b1 : n6206_o;
  assign n6208_o = n1909_o[80];
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6209_o = n6095_o ? n6208_o : n6134_o;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6211_o = n6095_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6213_o = n6095_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6215_o = n6095_o ? 1'b0 : n6180_o;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6217_o = n6095_o ? 1'b0 : n6182_o;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6219_o = n6095_o ? 2'b00 : n6184_o;
  /* TG68KdotC_Kernel.vhd:2781:41  */
  assign n6220_o = n6095_o ? n2180_o : n6185_o;
  /* TG68KdotC_Kernel.vhd:2823:50  */
  assign n6221_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2823:62  */
  assign n6223_o = n6221_o != 2'b11;
  /* TG68KdotC_Kernel.vhd:2824:52  */
  assign n6224_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:2824:55  */
  assign n6225_o = ~n6224_o;
  /* TG68KdotC_Kernel.vhd:2824:70  */
  assign n6226_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2824:82  */
  assign n6228_o = n6226_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2824:60  */
  assign n6229_o = n6228_o & n6225_o;
  /* TG68KdotC_Kernel.vhd:2824:101  */
  assign n6230_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2824:113  */
  assign n6232_o = n6230_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2824:131  */
  assign n6233_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:2824:143  */
  assign n6235_o = n6233_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2824:122  */
  assign n6236_o = n6232_o | n6235_o;
  /* TG68KdotC_Kernel.vhd:2824:90  */
  assign n6237_o = n6236_o & n6229_o;
  /* TG68KdotC_Kernel.vhd:2825:51  */
  assign n6238_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:2825:69  */
  assign n6239_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2825:81  */
  assign n6241_o = n6239_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:2825:59  */
  assign n6242_o = n6241_o & n6238_o;
  /* TG68KdotC_Kernel.vhd:2825:99  */
  assign n6243_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2825:111  */
  assign n6245_o = n6243_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:2825:128  */
  assign n6246_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2825:140  */
  assign n6248_o = n6246_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2825:119  */
  assign n6249_o = n6245_o | n6248_o;
  /* TG68KdotC_Kernel.vhd:2825:88  */
  assign n6250_o = n6249_o & n6242_o;
  /* TG68KdotC_Kernel.vhd:2824:151  */
  assign n6251_o = n6237_o | n6250_o;
  /* TG68KdotC_Kernel.vhd:2823:69  */
  assign n6252_o = n6251_o & n6223_o;
  /* TG68KdotC_Kernel.vhd:2823:41  */
  assign n6256_o = n6252_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2823:41  */
  assign n6259_o = n6252_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2823:41  */
  assign n6262_o = n6252_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2823:41  */
  assign n6264_o = n6252_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6265_o = n6092_o ? n6186_o : n1921_o;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6266_o = n6092_o ? n6187_o : datatype;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6268_o = n6092_o ? n6189_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6270_o = n6092_o ? n6191_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6272_o = n6092_o ? n6193_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6273_o = n6092_o ? n6194_o : n2154_o;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6274_o = n6092_o ? n6196_o : n6256_o;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6275_o = n6092_o ? n6198_o : n6259_o;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6277_o = n6092_o ? 1'b0 : n6262_o;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6279_o = n6092_o ? n6201_o : 1'b0;
  assign n6280_o = n1909_o[44];
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6281_o = n6092_o ? n6203_o : n6280_o;
  assign n6282_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6283_o = n6092_o ? n6205_o : n6282_o;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6285_o = n6095_o & n6092_o;
  assign n6286_o = n1909_o[80];
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6287_o = n6092_o ? n6209_o : n6286_o;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6289_o = n6092_o ? n6211_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6291_o = n6092_o ? 1'b0 : n6264_o;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6293_o = n6092_o ? n6213_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6295_o = n6092_o ? n6215_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6297_o = n6092_o ? n6217_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6299_o = n6092_o ? n6219_o : 2'b00;
  /* TG68KdotC_Kernel.vhd:2780:33  */
  assign n6300_o = n6092_o ? n6220_o : n2180_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6301_o = n6020_o ? n6067_o : n6265_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6302_o = n6020_o ? datatype : n6266_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6303_o = n6068_o & n6020_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6305_o = n6020_o ? n6070_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6307_o = n6020_o ? 1'b0 : n6268_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6308_o = n6020_o ? n6073_o : n6270_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6309_o = n6020_o ? n6075_o : n6272_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6310_o = n6020_o ? n2154_o : n6273_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6311_o = n6020_o ? n6078_o : n6274_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6312_o = n6020_o ? n6081_o : n6275_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6314_o = n6020_o ? n6084_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6316_o = n6020_o ? 1'b0 : n6277_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6318_o = n6020_o ? 1'b0 : n6279_o;
  assign n6319_o = n1909_o[44];
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6320_o = n6020_o ? n6319_o : n6281_o;
  assign n6321_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6322_o = n6020_o ? n6321_o : n6283_o;
  assign n6323_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6324_o = n6020_o ? n6323_o : n6207_o;
  assign n6325_o = n1909_o[80];
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6326_o = n6020_o ? n6325_o : n6287_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6328_o = n6020_o ? 1'b0 : n6289_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6330_o = n6020_o ? 1'b0 : n6291_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6332_o = n6020_o ? 1'b0 : n6293_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6334_o = n6020_o ? 1'b0 : n6295_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6335_o = n6020_o ? n6086_o : n6297_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6337_o = n6020_o ? 2'b00 : n6299_o;
  /* TG68KdotC_Kernel.vhd:2757:33  */
  assign n6338_o = n6020_o ? n6051_o : n6300_o;
  /* TG68KdotC_Kernel.vhd:2756:25  */
  assign n6340_o = n2185_o == 4'b1000;
  /* TG68KdotC_Kernel.vhd:2836:42  */
  assign n6341_o = opcode[8:3];
  /* TG68KdotC_Kernel.vhd:2836:54  */
  assign n6343_o = n6341_o != 6'b000001;
  /* TG68KdotC_Kernel.vhd:2837:45  */
  assign n6344_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:2837:48  */
  assign n6345_o = ~n6344_o;
  /* TG68KdotC_Kernel.vhd:2837:62  */
  assign n6346_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2837:74  */
  assign n6348_o = n6346_o == 2'b11;
  /* TG68KdotC_Kernel.vhd:2837:53  */
  assign n6349_o = n6345_o | n6348_o;
  /* TG68KdotC_Kernel.vhd:2837:92  */
  assign n6350_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2837:104  */
  assign n6352_o = n6350_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2837:122  */
  assign n6353_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:2837:134  */
  assign n6355_o = n6353_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2837:113  */
  assign n6356_o = n6352_o | n6355_o;
  /* TG68KdotC_Kernel.vhd:2837:81  */
  assign n6357_o = n6356_o & n6349_o;
  /* TG68KdotC_Kernel.vhd:2838:43  */
  assign n6358_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:2838:62  */
  assign n6359_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2838:74  */
  assign n6361_o = n6359_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:2838:91  */
  assign n6362_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2838:103  */
  assign n6364_o = n6362_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2838:82  */
  assign n6365_o = n6361_o | n6364_o;
  /* TG68KdotC_Kernel.vhd:2838:51  */
  assign n6366_o = n6365_o & n6358_o;
  /* TG68KdotC_Kernel.vhd:2837:142  */
  assign n6367_o = n6357_o | n6366_o;
  /* TG68KdotC_Kernel.vhd:2836:65  */
  assign n6368_o = n6367_o & n6343_o;
  /* TG68KdotC_Kernel.vhd:2841:50  */
  assign n6370_o = opcode[14];
  /* TG68KdotC_Kernel.vhd:2841:54  */
  assign n6371_o = ~n6370_o;
  assign n6373_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6374_o = n6448_o ? 1'b1 : n6373_o;
  /* TG68KdotC_Kernel.vhd:2844:50  */
  assign n6375_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2844:62  */
  assign n6377_o = n6375_o == 2'b11;
  /* TG68KdotC_Kernel.vhd:2845:58  */
  assign n6378_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:2845:61  */
  assign n6379_o = ~n6378_o;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6381_o = n6423_o ? 2'b01 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2850:58  */
  assign n6383_o = opcode[3];
  /* TG68KdotC_Kernel.vhd:2850:49  */
  assign n6386_o = n6383_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2854:49  */
  assign n6390_o = setexecopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2854:49  */
  assign n6393_o = setexecopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2859:58  */
  assign n6394_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:2859:76  */
  assign n6395_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2859:88  */
  assign n6397_o = n6395_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2859:66  */
  assign n6398_o = n6397_o & n6394_o;
  /* TG68KdotC_Kernel.vhd:2859:49  */
  assign n6401_o = n6398_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2859:49  */
  assign n6404_o = n6398_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2844:41  */
  assign n6405_o = n6379_o & n6377_o;
  /* TG68KdotC_Kernel.vhd:2844:41  */
  assign n6407_o = n6377_o ? n6386_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2844:41  */
  assign n6410_o = n6377_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2844:41  */
  assign n6412_o = n6377_o ? n6390_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2844:41  */
  assign n6414_o = n6377_o ? n6393_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2844:41  */
  assign n6416_o = n6377_o ? 1'b0 : n6401_o;
  /* TG68KdotC_Kernel.vhd:2844:41  */
  assign n6418_o = n6377_o ? 1'b0 : n6404_o;
  assign n6419_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6420_o = n6446_o ? 1'b1 : n6419_o;
  /* TG68KdotC_Kernel.vhd:2844:41  */
  assign n6422_o = n6377_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6423_o = n6405_o & n6368_o;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6425_o = n6368_o ? n6407_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6427_o = n6368_o ? n6410_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6429_o = n6368_o ? n6412_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6431_o = n6368_o ? n6414_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6434_o = n6368_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6437_o = n6368_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6440_o = n6368_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6442_o = n6368_o ? n6416_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6444_o = n6368_o ? n6418_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6446_o = n6377_o & n6368_o;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6448_o = n6371_o & n6368_o;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6450_o = n6368_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2836:33  */
  assign n6452_o = n6368_o ? n6422_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2835:25  */
  assign n6454_o = n2185_o == 4'b1001;
  /* TG68KdotC_Kernel.vhd:2835:36  */
  assign n6456_o = n2185_o == 4'b1101;
  /* TG68KdotC_Kernel.vhd:2835:36  */
  assign n6457_o = n6454_o | n6456_o;
  /* TG68KdotC_Kernel.vhd:2871:25  */
  assign n6459_o = n2185_o == 4'b1010;
  /* TG68KdotC_Kernel.vhd:2876:42  */
  assign n6460_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2876:54  */
  assign n6462_o = n6460_o == 2'b11;
  /* TG68KdotC_Kernel.vhd:2877:50  */
  assign n6463_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2877:62  */
  assign n6465_o = n6463_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2877:80  */
  assign n6466_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:2877:92  */
  assign n6468_o = n6466_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2877:71  */
  assign n6469_o = n6465_o | n6468_o;
  /* TG68KdotC_Kernel.vhd:2879:58  */
  assign n6470_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:2879:61  */
  assign n6471_o = ~n6470_o;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6474_o = n6638_o ? 2'b01 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2879:49  */
  assign n6476_o = n6471_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2886:66  */
  assign n6478_o = opcode[3];
  /* TG68KdotC_Kernel.vhd:2886:57  */
  assign n6481_o = n6478_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2884:49  */
  assign n6483_o = setexecopc ? n6481_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2884:49  */
  assign n6486_o = setexecopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2884:49  */
  assign n6489_o = setexecopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2884:49  */
  assign n6492_o = setexecopc ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2877:41  */
  assign n6494_o = n6471_o & n6469_o;
  /* TG68KdotC_Kernel.vhd:2877:41  */
  assign n6496_o = n6469_o ? n6483_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2877:41  */
  assign n6498_o = n6469_o ? n6486_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2877:41  */
  assign n6500_o = n6469_o ? n6489_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2877:41  */
  assign n6502_o = n6469_o ? n6492_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2877:41  */
  assign n6505_o = n6469_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2877:41  */
  assign n6508_o = n6469_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2877:41  */
  assign n6511_o = n6469_o ? 1'b1 : 1'b0;
  assign n6512_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2877:41  */
  assign n6513_o = n6469_o ? 1'b1 : n6512_o;
  /* TG68KdotC_Kernel.vhd:2877:41  */
  assign n6515_o = n6469_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2877:41  */
  assign n6517_o = n6469_o ? n6476_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2898:50  */
  assign n6518_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:2899:58  */
  assign n6519_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2899:70  */
  assign n6521_o = n6519_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:2903:74  */
  assign n6523_o = opcode[2:0];
  /* TG68KdotC_Kernel.vhd:2903:86  */
  assign n6525_o = n6523_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6527_o = n6627_o ? 1'b1 : n2168_o;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6531_o = n6617_o ? 2'b10 : n2026_o;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6532_o = n6622_o ? 1'b1 : n2007_o;
  assign n6533_o = n2162_o[0];
  assign n6534_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n6535_o = n2037_o ? n6533_o : n6534_o;
  /* TG68KdotC_Kernel.vhd:2902:57  */
  assign n6536_o = decodeopc ? 1'b1 : n6535_o;
  /* TG68KdotC_Kernel.vhd:2902:57  */
  assign n6537_o = n6525_o & decodeopc;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6539_o = n6637_o ? 7'b0100010 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2914:66  */
  assign n6542_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2914:78  */
  assign n6544_o = n6542_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:2914:95  */
  assign n6545_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2914:107  */
  assign n6547_o = n6545_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2914:86  */
  assign n6548_o = n6544_o | n6547_o;
  /* TG68KdotC_Kernel.vhd:2914:57  */
  assign n6552_o = n6548_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2914:57  */
  assign n6555_o = n6548_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2914:57  */
  assign n6558_o = n6548_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2914:57  */
  assign n6561_o = n6548_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2914:57  */
  assign n6563_o = n6548_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2899:49  */
  assign n6564_o = decodeopc & n6521_o;
  /* TG68KdotC_Kernel.vhd:2899:49  */
  assign n6566_o = n6521_o ? 1'b0 : n6552_o;
  /* TG68KdotC_Kernel.vhd:2899:49  */
  assign n6568_o = n6521_o ? 1'b0 : n6555_o;
  /* TG68KdotC_Kernel.vhd:2899:49  */
  assign n6570_o = n6521_o ? 1'b1 : n6558_o;
  /* TG68KdotC_Kernel.vhd:2899:49  */
  assign n6572_o = n6521_o ? 1'b0 : n6561_o;
  /* TG68KdotC_Kernel.vhd:2899:49  */
  assign n6573_o = decodeopc & n6521_o;
  assign n6574_o = n2162_o[0];
  assign n6575_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n6576_o = n2037_o ? n6574_o : n6575_o;
  /* TG68KdotC_Kernel.vhd:2899:49  */
  assign n6577_o = n6521_o ? n6536_o : n6576_o;
  /* TG68KdotC_Kernel.vhd:2899:49  */
  assign n6578_o = n6537_o & n6521_o;
  assign n6579_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2899:49  */
  assign n6580_o = n6521_o ? 1'b1 : n6579_o;
  /* TG68KdotC_Kernel.vhd:2899:49  */
  assign n6582_o = n6521_o ? 1'b0 : n6563_o;
  /* TG68KdotC_Kernel.vhd:2899:49  */
  assign n6584_o = n6521_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2899:49  */
  assign n6586_o = n6521_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2899:49  */
  assign n6587_o = decodeopc & n6521_o;
  /* TG68KdotC_Kernel.vhd:2924:58  */
  assign n6588_o = opcode[8:3];
  /* TG68KdotC_Kernel.vhd:2924:70  */
  assign n6590_o = n6588_o != 6'b000001;
  /* TG68KdotC_Kernel.vhd:2925:59  */
  assign n6591_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2925:71  */
  assign n6593_o = n6591_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2925:89  */
  assign n6594_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:2925:101  */
  assign n6596_o = n6594_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2925:80  */
  assign n6597_o = n6593_o | n6596_o;
  /* TG68KdotC_Kernel.vhd:2924:81  */
  assign n6598_o = n6597_o & n6590_o;
  /* TG68KdotC_Kernel.vhd:2924:49  */
  assign n6603_o = n6598_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2924:49  */
  assign n6606_o = n6598_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2924:49  */
  assign n6609_o = n6598_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2924:49  */
  assign n6612_o = n6598_o ? 1'b1 : 1'b0;
  assign n6613_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:2924:49  */
  assign n6614_o = n6598_o ? 1'b1 : n6613_o;
  /* TG68KdotC_Kernel.vhd:2924:49  */
  assign n6616_o = n6598_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6617_o = n6564_o & n6518_o;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6618_o = n6518_o ? n6566_o : n6603_o;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6619_o = n6518_o ? n6568_o : n6606_o;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6620_o = n6518_o ? n6570_o : n6609_o;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6621_o = n6518_o ? n6572_o : n6612_o;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6622_o = n6573_o & n6518_o;
  assign n6623_o = n2162_o[0];
  assign n6624_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n6625_o = n2037_o ? n6623_o : n6624_o;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6626_o = n6518_o ? n6577_o : n6625_o;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6627_o = n6578_o & n6518_o;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6628_o = n6518_o ? n6580_o : n6614_o;
  assign n6629_o = {n6584_o, n6582_o};
  assign n6630_o = n6629_o[0];
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6632_o = n6518_o ? n6630_o : 1'b0;
  assign n6633_o = n6629_o[1];
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6634_o = n6518_o ? n6633_o : n6616_o;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6636_o = n6518_o ? n6586_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2898:41  */
  assign n6637_o = n6587_o & n6518_o;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6638_o = n6494_o & n6462_o;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6639_o = n6462_o ? n2026_o : n6531_o;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6641_o = n6462_o ? n6496_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6643_o = n6462_o ? n6498_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6645_o = n6462_o ? n6500_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6647_o = n6462_o ? n6502_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6648_o = n6462_o ? n6505_o : n6618_o;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6649_o = n6462_o ? n6508_o : n6619_o;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6650_o = n6462_o ? n6511_o : n6620_o;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6652_o = n6462_o ? 1'b0 : n6621_o;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6653_o = n6462_o ? n2007_o : n6532_o;
  assign n6654_o = n2162_o[0];
  assign n6655_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n6656_o = n2037_o ? n6654_o : n6655_o;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6657_o = n6462_o ? n6656_o : n6626_o;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6658_o = n6462_o ? n2168_o : n6527_o;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6659_o = n6462_o ? n6513_o : n6628_o;
  assign n6660_o = {n6634_o, n6632_o};
  assign n6661_o = n6660_o[0];
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6663_o = n6462_o ? 1'b0 : n6661_o;
  assign n6664_o = n6660_o[1];
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6665_o = n6462_o ? n6515_o : n6664_o;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6667_o = n6462_o ? n6517_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6669_o = n6462_o ? 1'b0 : n6636_o;
  /* TG68KdotC_Kernel.vhd:2876:33  */
  assign n6670_o = n6462_o ? n2180_o : n6539_o;
  /* TG68KdotC_Kernel.vhd:2875:25  */
  assign n6672_o = n2185_o == 4'b1011;
  /* TG68KdotC_Kernel.vhd:2939:42  */
  assign n6673_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2939:54  */
  assign n6675_o = n6673_o == 2'b11;
  /* TG68KdotC_Kernel.vhd:2941:50  */
  assign n6676_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2941:62  */
  assign n6678_o = n6676_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2940:56  */
  assign n6680_o = n6678_o & 1'b1;
  /* TG68KdotC_Kernel.vhd:2941:81  */
  assign n6681_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2941:93  */
  assign n6683_o = n6681_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2941:111  */
  assign n6684_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:2941:123  */
  assign n6686_o = n6684_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2941:102  */
  assign n6687_o = n6683_o | n6686_o;
  /* TG68KdotC_Kernel.vhd:2941:70  */
  assign n6688_o = n6687_o & n6680_o;
  /* TG68KdotC_Kernel.vhd:2942:58  */
  assign n6689_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2942:70  */
  assign n6691_o = n6689_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2942:49  */
  assign n6694_o = n6691_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2945:64  */
  assign n6696_o = micro_state == 7'b0000000;
  /* TG68KdotC_Kernel.vhd:2945:70  */
  assign n6697_o = nextpass & n6696_o;
  /* TG68KdotC_Kernel.vhd:2945:98  */
  assign n6698_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2945:110  */
  assign n6700_o = n6698_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2945:116  */
  assign n6701_o = decodeopc & n6700_o;
  /* TG68KdotC_Kernel.vhd:2945:88  */
  assign n6702_o = n6697_o | n6701_o;
  /* TG68KdotC_Kernel.vhd:2940:41  */
  assign n6705_o = n6724_o ? 2'b01 : n2026_o;
  assign n6706_o = n1909_o[24];
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n6707_o = n6916_o ? 1'b1 : n6706_o;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n6709_o = n6931_o ? 7'b1010101 : n2180_o;
  /* TG68KdotC_Kernel.vhd:2958:77  */
  assign n6711_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2958:89  */
  assign n6713_o = n6711_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2958:95  */
  assign n6714_o = decodeopc & n6713_o;
  /* TG68KdotC_Kernel.vhd:2958:67  */
  assign n6715_o = nextpass | n6714_o;
  /* TG68KdotC_Kernel.vhd:2958:49  */
  assign n6718_o = n6715_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2962:49  */
  assign n6721_o = setexecopc ? 2'b10 : 2'b01;
  /* TG68KdotC_Kernel.vhd:2940:41  */
  assign n6723_o = n6688_o ? n6721_o : n1921_o;
  /* TG68KdotC_Kernel.vhd:2940:41  */
  assign n6724_o = n6702_o & n6688_o;
  /* TG68KdotC_Kernel.vhd:2940:41  */
  assign n6726_o = n6688_o ? n6694_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2940:41  */
  assign n6729_o = n6688_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2940:41  */
  assign n6731_o = n6688_o ? n6718_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2940:41  */
  assign n6734_o = n6688_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2940:41  */
  assign n6737_o = n6688_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2940:41  */
  assign n6740_o = n6688_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2940:41  */
  assign n6742_o = n6702_o & n6688_o;
  /* TG68KdotC_Kernel.vhd:2940:41  */
  assign n6744_o = n6688_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2940:41  */
  assign n6745_o = n6702_o & n6688_o;
  /* TG68KdotC_Kernel.vhd:2969:45  */
  assign n6746_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:2969:63  */
  assign n6747_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2969:75  */
  assign n6749_o = n6747_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2969:53  */
  assign n6750_o = n6749_o & n6746_o;
  /* TG68KdotC_Kernel.vhd:2970:50  */
  assign n6751_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2970:62  */
  assign n6753_o = n6751_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2975:58  */
  assign n6756_o = opcode[7:4];
  /* TG68KdotC_Kernel.vhd:2975:70  */
  assign n6758_o = n6756_o == 4'b0100;
  /* TG68KdotC_Kernel.vhd:2975:87  */
  assign n6759_o = opcode[7:3];
  /* TG68KdotC_Kernel.vhd:2975:99  */
  assign n6761_o = n6759_o == 5'b10001;
  /* TG68KdotC_Kernel.vhd:2975:78  */
  assign n6762_o = n6758_o | n6761_o;
  /* TG68KdotC_Kernel.vhd:2980:66  */
  assign n6766_o = opcode[6];
  /* TG68KdotC_Kernel.vhd:2980:84  */
  assign n6767_o = opcode[3];
  /* TG68KdotC_Kernel.vhd:2980:74  */
  assign n6768_o = n6767_o & n6766_o;
  /* TG68KdotC_Kernel.vhd:2980:57  */
  assign n6771_o = n6768_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2980:57  */
  assign n6774_o = n6768_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2975:49  */
  assign n6776_o = n6782_o ? 2'b01 : n2026_o;
  /* TG68KdotC_Kernel.vhd:2984:57  */
  assign n6779_o = decodeopc ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2975:49  */
  assign n6781_o = n6762_o ? 2'b10 : n1921_o;
  /* TG68KdotC_Kernel.vhd:2975:49  */
  assign n6782_o = decodeopc & n6762_o;
  /* TG68KdotC_Kernel.vhd:2975:49  */
  assign n6784_o = n6762_o ? n6771_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2975:49  */
  assign n6786_o = n6762_o ? n6774_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2975:49  */
  assign n6788_o = n6762_o ? n6779_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2975:49  */
  assign n6791_o = n6762_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2975:49  */
  assign n6794_o = n6762_o ? 1'b0 : 1'b1;
  assign n6795_o = n1909_o[34];
  /* TG68KdotC_Kernel.vhd:2975:49  */
  assign n6796_o = n6762_o ? 1'b1 : n6795_o;
  assign n6797_o = n1909_o[61];
  /* TG68KdotC_Kernel.vhd:2975:49  */
  assign n6798_o = n6762_o ? 1'b1 : n6797_o;
  assign n6799_o = n1909_o[85];
  /* TG68KdotC_Kernel.vhd:2975:49  */
  assign n6800_o = n6762_o ? 1'b1 : n6799_o;
  /* TG68KdotC_Kernel.vhd:2970:41  */
  assign n6801_o = n6753_o ? n1921_o : n6781_o;
  /* TG68KdotC_Kernel.vhd:2970:41  */
  assign n6802_o = n6753_o ? n2026_o : n6776_o;
  /* TG68KdotC_Kernel.vhd:2970:41  */
  assign n6804_o = n6753_o ? 1'b0 : n6784_o;
  /* TG68KdotC_Kernel.vhd:2970:41  */
  assign n6806_o = n6753_o ? 1'b0 : n6786_o;
  /* TG68KdotC_Kernel.vhd:2970:41  */
  assign n6808_o = n6753_o ? 1'b0 : n6788_o;
  /* TG68KdotC_Kernel.vhd:2970:41  */
  assign n6810_o = n6753_o ? 1'b0 : n6791_o;
  /* TG68KdotC_Kernel.vhd:2970:41  */
  assign n6812_o = n6753_o ? 1'b0 : n6794_o;
  /* TG68KdotC_Kernel.vhd:2970:41  */
  assign n6815_o = n6753_o ? 1'b1 : 1'b0;
  assign n6816_o = n1909_o[34];
  /* TG68KdotC_Kernel.vhd:2970:41  */
  assign n6817_o = n6753_o ? n6816_o : n6796_o;
  assign n6818_o = n1909_o[61];
  /* TG68KdotC_Kernel.vhd:2970:41  */
  assign n6819_o = n6753_o ? n6818_o : n6798_o;
  assign n6820_o = n1909_o[85];
  /* TG68KdotC_Kernel.vhd:2970:41  */
  assign n6821_o = n6753_o ? n6820_o : n6800_o;
  /* TG68KdotC_Kernel.vhd:2970:41  */
  assign n6823_o = n6753_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2970:41  */
  assign n6825_o = n6753_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2995:50  */
  assign n6826_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:2995:62  */
  assign n6828_o = n6826_o != 2'b11;
  /* TG68KdotC_Kernel.vhd:2996:52  */
  assign n6829_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:2996:55  */
  assign n6830_o = ~n6829_o;
  /* TG68KdotC_Kernel.vhd:2996:70  */
  assign n6831_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2996:82  */
  assign n6833_o = n6831_o != 3'b001;
  /* TG68KdotC_Kernel.vhd:2996:60  */
  assign n6834_o = n6833_o & n6830_o;
  /* TG68KdotC_Kernel.vhd:2996:101  */
  assign n6835_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:2996:113  */
  assign n6837_o = n6835_o != 4'b1111;
  /* TG68KdotC_Kernel.vhd:2996:131  */
  assign n6838_o = opcode[1:0];
  /* TG68KdotC_Kernel.vhd:2996:143  */
  assign n6840_o = n6838_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2996:122  */
  assign n6841_o = n6837_o | n6840_o;
  /* TG68KdotC_Kernel.vhd:2996:90  */
  assign n6842_o = n6841_o & n6834_o;
  /* TG68KdotC_Kernel.vhd:2997:51  */
  assign n6843_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:2997:69  */
  assign n6844_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:2997:81  */
  assign n6846_o = n6844_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:2997:59  */
  assign n6847_o = n6846_o & n6843_o;
  /* TG68KdotC_Kernel.vhd:2997:99  */
  assign n6848_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:2997:111  */
  assign n6850_o = n6848_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:2997:128  */
  assign n6851_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:2997:140  */
  assign n6853_o = n6851_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:2997:119  */
  assign n6854_o = n6850_o | n6853_o;
  /* TG68KdotC_Kernel.vhd:2997:88  */
  assign n6855_o = n6854_o & n6847_o;
  /* TG68KdotC_Kernel.vhd:2996:151  */
  assign n6856_o = n6842_o | n6855_o;
  /* TG68KdotC_Kernel.vhd:2995:69  */
  assign n6857_o = n6856_o & n6828_o;
  /* TG68KdotC_Kernel.vhd:2995:41  */
  assign n6861_o = n6857_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2995:41  */
  assign n6864_o = n6857_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:2995:41  */
  assign n6867_o = n6857_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2995:41  */
  assign n6869_o = n6857_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n6870_o = n6750_o ? n6801_o : n1921_o;
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n6871_o = n6750_o ? n6802_o : n2026_o;
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n6873_o = n6750_o ? n6804_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n6875_o = n6750_o ? n6806_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n6877_o = n6750_o ? n6808_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n6878_o = n6750_o ? n6810_o : n6861_o;
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n6879_o = n6750_o ? n6812_o : n6864_o;
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n6881_o = n6750_o ? 1'b0 : n6867_o;
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n6883_o = n6750_o ? n6815_o : 1'b0;
  assign n6884_o = n1909_o[34];
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n6885_o = n6750_o ? n6817_o : n6884_o;
  assign n6886_o = n1909_o[61];
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n6887_o = n6750_o ? n6819_o : n6886_o;
  assign n6888_o = n1909_o[85];
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n6889_o = n6750_o ? n6821_o : n6888_o;
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n6891_o = n6750_o ? n6823_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n6893_o = n6750_o ? 1'b0 : n6869_o;
  /* TG68KdotC_Kernel.vhd:2969:33  */
  assign n6895_o = n6750_o ? n6825_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n6896_o = n6675_o ? n6723_o : n6870_o;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n6897_o = n6675_o ? n6705_o : n6871_o;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n6899_o = n6675_o ? n6726_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n6901_o = n6675_o ? 1'b0 : n6873_o;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n6903_o = n6675_o ? n6729_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n6905_o = n6675_o ? 1'b0 : n6875_o;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n6906_o = n6675_o ? n6731_o : n6877_o;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n6907_o = n6675_o ? n6734_o : n6878_o;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n6908_o = n6675_o ? n6737_o : n6879_o;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n6910_o = n6675_o ? n6740_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n6912_o = n6675_o ? 1'b0 : n6881_o;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n6914_o = n6675_o ? 1'b0 : n6883_o;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n6916_o = n6742_o & n6675_o;
  assign n6917_o = n1909_o[34];
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n6918_o = n6675_o ? n6917_o : n6885_o;
  assign n6919_o = n1909_o[61];
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n6920_o = n6675_o ? n6919_o : n6887_o;
  assign n6921_o = n1909_o[85];
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n6922_o = n6675_o ? n6921_o : n6889_o;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n6924_o = n6675_o ? 1'b0 : n6891_o;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n6926_o = n6675_o ? 1'b0 : n6893_o;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n6928_o = n6675_o ? 1'b0 : n6895_o;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n6930_o = n6675_o ? n6744_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:2939:33  */
  assign n6931_o = n6745_o & n6675_o;
  /* TG68KdotC_Kernel.vhd:2938:25  */
  assign n6933_o = n2185_o == 4'b1100;
  /* TG68KdotC_Kernel.vhd:3008:42  */
  assign n6934_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:3008:54  */
  assign n6936_o = n6934_o == 2'b11;
  /* TG68KdotC_Kernel.vhd:3009:50  */
  assign n6937_o = opcode[11];
  /* TG68KdotC_Kernel.vhd:3009:54  */
  assign n6938_o = ~n6937_o;
  /* TG68KdotC_Kernel.vhd:3010:54  */
  assign n6939_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:3010:66  */
  assign n6941_o = n6939_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:3010:84  */
  assign n6942_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:3010:96  */
  assign n6944_o = n6942_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:3010:113  */
  assign n6945_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:3010:125  */
  assign n6947_o = n6945_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:3010:104  */
  assign n6948_o = n6944_o | n6947_o;
  /* TG68KdotC_Kernel.vhd:3010:73  */
  assign n6949_o = n6948_o & n6941_o;
  /* TG68KdotC_Kernel.vhd:3018:79  */
  assign n6951_o = opcode[10:9];
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n6954_o = n7265_o ? 2'b01 : n1921_o;
  /* TG68KdotC_Kernel.vhd:3010:44  */
  assign n6957_o = n6949_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n6958_o = n7282_o ? n6951_o : n1900_o;
  /* TG68KdotC_Kernel.vhd:3010:44  */
  assign n6961_o = n6949_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3010:44  */
  assign n6964_o = n6949_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3010:44  */
  assign n6967_o = n6949_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3010:44  */
  assign n6969_o = n6949_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3010:44  */
  assign n6971_o = n6949_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3026:70  */
  assign n6972_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:3026:73  */
  assign n6973_o = ~n6972_o;
  /* TG68KdotC_Kernel.vhd:3026:78  */
  assign n6975_o = 1'b1 & n6973_o;
  /* TG68KdotC_Kernel.vhd:3026:63  */
  assign n6977_o = 1'b0 | n6975_o;
  /* TG68KdotC_Kernel.vhd:3027:60  */
  assign n6978_o = opcode[10:9];
  /* TG68KdotC_Kernel.vhd:3027:73  */
  assign n6980_o = n6978_o == 2'b11;
  /* TG68KdotC_Kernel.vhd:3027:88  */
  assign n6981_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3027:101  */
  assign n6983_o = n6981_o == 3'b010;
  /* TG68KdotC_Kernel.vhd:3027:79  */
  assign n6984_o = n6980_o | n6983_o;
  /* TG68KdotC_Kernel.vhd:3027:117  */
  assign n6985_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3027:130  */
  assign n6987_o = n6985_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:3027:108  */
  assign n6988_o = n6984_o | n6987_o;
  /* TG68KdotC_Kernel.vhd:3028:59  */
  assign n6989_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:3028:71  */
  assign n6991_o = n6989_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:3028:87  */
  assign n6992_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:3028:99  */
  assign n6994_o = n6992_o == 3'b011;
  /* TG68KdotC_Kernel.vhd:3028:78  */
  assign n6995_o = n6991_o | n6994_o;
  /* TG68KdotC_Kernel.vhd:3028:115  */
  assign n6996_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:3028:127  */
  assign n6998_o = n6996_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:3028:106  */
  assign n6999_o = n6995_o | n6998_o;
  /* TG68KdotC_Kernel.vhd:3028:144  */
  assign n7000_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:3028:156  */
  assign n7002_o = n7000_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:3028:173  */
  assign n7003_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:3028:185  */
  assign n7005_o = n7003_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:3028:163  */
  assign n7006_o = n7005_o & n7002_o;
  /* TG68KdotC_Kernel.vhd:3028:134  */
  assign n7007_o = n6999_o | n7006_o;
  /* TG68KdotC_Kernel.vhd:3027:138  */
  assign n7008_o = n7007_o & n6988_o;
  /* TG68KdotC_Kernel.vhd:3026:94  */
  assign n7009_o = n6977_o | n7008_o;
  /* TG68KdotC_Kernel.vhd:3029:60  */
  assign n7010_o = opcode[10:9];
  /* TG68KdotC_Kernel.vhd:3029:73  */
  assign n7012_o = n7010_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:3029:88  */
  assign n7013_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3029:101  */
  assign n7015_o = n7013_o == 3'b011;
  /* TG68KdotC_Kernel.vhd:3029:79  */
  assign n7016_o = n7012_o | n7015_o;
  /* TG68KdotC_Kernel.vhd:3029:117  */
  assign n7017_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3029:130  */
  assign n7019_o = n7017_o == 3'b101;
  /* TG68KdotC_Kernel.vhd:3029:108  */
  assign n7020_o = n7016_o | n7019_o;
  /* TG68KdotC_Kernel.vhd:3030:59  */
  assign n7021_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:3030:71  */
  assign n7023_o = n7021_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:3030:87  */
  assign n7024_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:3030:99  */
  assign n7026_o = n7024_o == 3'b011;
  /* TG68KdotC_Kernel.vhd:3030:78  */
  assign n7027_o = n7023_o | n7026_o;
  /* TG68KdotC_Kernel.vhd:3030:115  */
  assign n7028_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:3030:127  */
  assign n7030_o = n7028_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:3030:106  */
  assign n7031_o = n7027_o | n7030_o;
  /* TG68KdotC_Kernel.vhd:3030:143  */
  assign n7032_o = opcode[5:2];
  /* TG68KdotC_Kernel.vhd:3030:155  */
  assign n7034_o = n7032_o == 4'b1111;
  /* TG68KdotC_Kernel.vhd:3030:134  */
  assign n7035_o = n7031_o | n7034_o;
  /* TG68KdotC_Kernel.vhd:3029:138  */
  assign n7036_o = n7035_o & n7020_o;
  /* TG68KdotC_Kernel.vhd:3028:195  */
  assign n7037_o = n7009_o | n7036_o;
  assign n7040_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:3034:57  */
  assign n7041_o = decodeopc ? 1'b1 : n7040_o;
  assign n7042_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:3034:57  */
  assign n7043_o = decodeopc ? 1'b1 : n7042_o;
  /* TG68KdotC_Kernel.vhd:3034:57  */
  assign n7045_o = decodeopc ? 7'b0000001 : n2180_o;
  /* TG68KdotC_Kernel.vhd:3041:66  */
  assign n7047_o = opcode[10];
  /* TG68KdotC_Kernel.vhd:3041:84  */
  assign n7048_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:3041:87  */
  assign n7049_o = ~n7048_o;
  /* TG68KdotC_Kernel.vhd:3041:75  */
  assign n7050_o = n7047_o | n7049_o;
  /* TG68KdotC_Kernel.vhd:3041:57  */
  assign n7053_o = n7050_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3044:66  */
  assign n7054_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3044:79  */
  assign n7056_o = n7054_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:3044:57  */
  assign n7059_o = n7056_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3047:66  */
  assign n7060_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3047:79  */
  assign n7062_o = n7060_o == 3'b010;
  /* TG68KdotC_Kernel.vhd:3047:95  */
  assign n7063_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3047:108  */
  assign n7065_o = n7063_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:3047:86  */
  assign n7066_o = n7062_o | n7065_o;
  /* TG68KdotC_Kernel.vhd:3047:124  */
  assign n7067_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3047:137  */
  assign n7069_o = n7067_o == 3'b110;
  /* TG68KdotC_Kernel.vhd:3047:115  */
  assign n7070_o = n7066_o | n7069_o;
  /* TG68KdotC_Kernel.vhd:3047:153  */
  assign n7071_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3047:166  */
  assign n7073_o = n7071_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:3047:144  */
  assign n7074_o = n7070_o | n7073_o;
  /* TG68KdotC_Kernel.vhd:3047:57  */
  assign n7077_o = n7074_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3051:66  */
  assign n7078_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3051:79  */
  assign n7080_o = n7078_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:3051:95  */
  assign n7081_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3051:108  */
  assign n7083_o = n7081_o == 3'b011;
  /* TG68KdotC_Kernel.vhd:3051:86  */
  assign n7084_o = n7080_o | n7083_o;
  /* TG68KdotC_Kernel.vhd:3051:124  */
  assign n7085_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3051:137  */
  assign n7087_o = n7085_o == 3'b101;
  /* TG68KdotC_Kernel.vhd:3051:115  */
  assign n7088_o = n7084_o | n7087_o;
  /* TG68KdotC_Kernel.vhd:3051:57  */
  assign n7091_o = n7088_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3054:66  */
  assign n7092_o = opcode[4:3];
  /* TG68KdotC_Kernel.vhd:3054:78  */
  assign n7094_o = n7092_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:3055:74  */
  assign n7095_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3055:87  */
  assign n7097_o = n7095_o != 3'b000;
  /* TG68KdotC_Kernel.vhd:3054:57  */
  assign n7099_o = n7119_o ? 1'b1 : n7091_o;
  /* TG68KdotC_Kernel.vhd:3058:72  */
  assign n7100_o = exec[42];
  /* TG68KdotC_Kernel.vhd:3054:57  */
  assign n7103_o = n7112_o ? 2'b01 : n2026_o;
  /* TG68KdotC_Kernel.vhd:3058:65  */
  assign n7106_o = n7100_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3058:65  */
  assign n7109_o = n7100_o ? 1'b1 : 1'b0;
  assign n7110_o = n1909_o[29];
  /* TG68KdotC_Kernel.vhd:3054:57  */
  assign n7111_o = n7118_o ? 1'b1 : n7110_o;
  /* TG68KdotC_Kernel.vhd:3054:57  */
  assign n7112_o = n7100_o & n7094_o;
  /* TG68KdotC_Kernel.vhd:3054:57  */
  assign n7114_o = n7094_o ? n7106_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3054:57  */
  assign n7116_o = n7094_o ? n7109_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3054:57  */
  assign n7118_o = n7100_o & n7094_o;
  /* TG68KdotC_Kernel.vhd:3054:57  */
  assign n7119_o = n7097_o & n7094_o;
  /* TG68KdotC_Kernel.vhd:3065:63  */
  assign n7120_o = set[62];
  /* TG68KdotC_Kernel.vhd:3065:57  */
  assign n7122_o = n7120_o ? 2'b01 : n7103_o;
  /* TG68KdotC_Kernel.vhd:3068:64  */
  assign n7123_o = exec[62];
  /* TG68KdotC_Kernel.vhd:3068:57  */
  assign n7127_o = n7123_o ? 2'b01 : n7122_o;
  /* TG68KdotC_Kernel.vhd:3068:57  */
  assign n7129_o = n7123_o ? 1'b1 : n7114_o;
  /* TG68KdotC_Kernel.vhd:3068:57  */
  assign n7131_o = n7123_o ? 1'b1 : n7116_o;
  /* TG68KdotC_Kernel.vhd:3068:57  */
  assign n7132_o = n7123_o ? 1'b1 : n7111_o;
  assign n7133_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:3068:57  */
  assign n7134_o = n7123_o ? 1'b1 : n7133_o;
  /* TG68KdotC_Kernel.vhd:3068:57  */
  assign n7136_o = n7123_o ? 7'b1010100 : n7045_o;
  /* TG68KdotC_Kernel.vhd:3077:74  */
  assign n7137_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3077:87  */
  assign n7139_o = n7137_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:3077:65  */
  assign n7142_o = n7139_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3077:65  */
  assign n7145_o = n7139_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3082:74  */
  assign n7146_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3082:87  */
  assign n7148_o = n7146_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:3082:103  */
  assign n7149_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3082:116  */
  assign n7151_o = n7149_o == 3'b011;
  /* TG68KdotC_Kernel.vhd:3082:94  */
  assign n7152_o = n7148_o | n7151_o;
  /* TG68KdotC_Kernel.vhd:3082:132  */
  assign n7153_o = opcode[10:8];
  /* TG68KdotC_Kernel.vhd:3082:145  */
  assign n7155_o = n7153_o == 3'b101;
  /* TG68KdotC_Kernel.vhd:3082:123  */
  assign n7156_o = n7152_o | n7155_o;
  /* TG68KdotC_Kernel.vhd:3076:57  */
  assign n7158_o = n7163_o ? 1'b1 : n7131_o;
  /* TG68KdotC_Kernel.vhd:3076:57  */
  assign n7160_o = setexecopc ? n7142_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3076:57  */
  assign n7162_o = setexecopc ? n7145_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3076:57  */
  assign n7163_o = n7156_o & setexecopc;
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7164_o = n7037_o ? n2026_o : n7127_o;
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7166_o = n7037_o ? 1'b0 : n7077_o;
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7169_o = n7037_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7171_o = n7037_o ? 1'b0 : n7160_o;
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7173_o = n7037_o ? 1'b0 : n7162_o;
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7175_o = n7037_o ? 1'b0 : n7129_o;
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7177_o = n7037_o ? 1'b0 : n7158_o;
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7180_o = n7037_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7183_o = n7037_o ? 1'b1 : 1'b0;
  assign n7184_o = n1909_o[29];
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7185_o = n7037_o ? n7184_o : n7132_o;
  assign n7186_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7187_o = n7037_o ? n7186_o : n7041_o;
  assign n7188_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7189_o = n7037_o ? n7188_o : n7134_o;
  assign n7190_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7191_o = n7037_o ? n7190_o : n7043_o;
  assign n7192_o = {n7053_o, 1'b1};
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7194_o = n7037_o ? 1'b0 : n7059_o;
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7196_o = n7037_o ? 1'b0 : n7099_o;
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7198_o = n7037_o ? 2'b00 : n7192_o;
  /* TG68KdotC_Kernel.vhd:3026:49  */
  assign n7199_o = n7037_o ? n2180_o : n7136_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7200_o = n6949_o & n6938_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7201_o = n6938_o ? n2026_o : n7164_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7202_o = n6938_o ? n6957_o : n7166_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7204_o = n6938_o ? 1'b0 : n7169_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7206_o = n6938_o ? 1'b0 : n7171_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7208_o = n6938_o ? 1'b0 : n7173_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7210_o = n6938_o ? 1'b0 : n7175_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7212_o = n6938_o ? 1'b0 : n7177_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7213_o = n6949_o & n6938_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7214_o = n6938_o ? n6961_o : n7180_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7215_o = n6938_o ? n6964_o : n7183_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7217_o = n6938_o ? n6967_o : 1'b0;
  assign n7218_o = n1909_o[29];
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7219_o = n6938_o ? n7218_o : n7185_o;
  assign n7220_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7221_o = n6938_o ? n7220_o : n7187_o;
  assign n7222_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7223_o = n6938_o ? n7222_o : n7189_o;
  assign n7224_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7225_o = n6938_o ? n7224_o : n7191_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7227_o = n6938_o ? n6969_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7228_o = n6938_o ? n6971_o : n7194_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7230_o = n6938_o ? 1'b0 : n7196_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7232_o = n6938_o ? 2'b00 : n7198_o;
  /* TG68KdotC_Kernel.vhd:3009:41  */
  assign n7233_o = n6938_o ? n2180_o : n7199_o;
  /* TG68KdotC_Kernel.vhd:3095:66  */
  assign n7237_o = opcode[5];
  /* TG68KdotC_Kernel.vhd:3100:98  */
  assign n7239_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:3101:74  */
  assign n7240_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:3101:87  */
  assign n7242_o = n7240_o == 3'b000;
  /* TG68KdotC_Kernel.vhd:3101:65  */
  assign n7245_o = n7242_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3094:49  */
  assign n7247_o = n7257_o ? 2'b01 : n2026_o;
  assign n7248_o = {n7245_o, n7239_o};
  assign n7249_o = n1904_o[3:0];
  assign n7250_o = n1905_o[3:0];
  /* TG68KdotC_Kernel.vhd:1495:17  */
  assign n7251_o = n1902_o ? n7249_o : n7250_o;
  /* TG68KdotC_Kernel.vhd:3095:57  */
  assign n7252_o = n7237_o ? n7251_o : n7248_o;
  assign n7253_o = n1909_o[24];
  /* TG68KdotC_Kernel.vhd:3094:49  */
  assign n7254_o = n7263_o ? 1'b1 : n7253_o;
  /* TG68KdotC_Kernel.vhd:3094:49  */
  assign n7256_o = n7264_o ? 7'b1010011 : n2180_o;
  /* TG68KdotC_Kernel.vhd:3094:49  */
  assign n7257_o = n7237_o & decodeopc;
  assign n7258_o = n1904_o[3:0];
  assign n7259_o = n1905_o[3:0];
  /* TG68KdotC_Kernel.vhd:1495:17  */
  assign n7260_o = n1902_o ? n7258_o : n7259_o;
  /* TG68KdotC_Kernel.vhd:3094:49  */
  assign n7261_o = decodeopc ? n7252_o : n7260_o;
  /* TG68KdotC_Kernel.vhd:3094:49  */
  assign n7263_o = n7237_o & decodeopc;
  /* TG68KdotC_Kernel.vhd:3094:49  */
  assign n7264_o = n7237_o & decodeopc;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7265_o = n7200_o & n6936_o;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7266_o = n6936_o ? n7201_o : n7247_o;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7269_o = n6936_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7271_o = n6936_o ? n7202_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7273_o = n6936_o ? n7204_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7275_o = n6936_o ? n7206_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7277_o = n6936_o ? n7208_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7279_o = n6936_o ? n7210_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7281_o = n6936_o ? n7212_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7282_o = n7213_o & n6936_o;
  assign n7283_o = n1904_o[3:0];
  assign n7284_o = n1905_o[3:0];
  /* TG68KdotC_Kernel.vhd:1495:17  */
  assign n7285_o = n1902_o ? n7283_o : n7284_o;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7286_o = n6936_o ? n7285_o : n7261_o;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7288_o = n6936_o ? n7214_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7290_o = n6936_o ? n7215_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7292_o = n6936_o ? n7217_o : 1'b0;
  assign n7293_o = n1909_o[24];
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7294_o = n6936_o ? n7293_o : n7254_o;
  assign n7295_o = n1909_o[29];
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7296_o = n6936_o ? n7219_o : n7295_o;
  assign n7297_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7298_o = n6936_o ? n7221_o : n7297_o;
  assign n7299_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7300_o = n6936_o ? n7223_o : n7299_o;
  assign n7301_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7302_o = n6936_o ? n7225_o : n7301_o;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7303_o = n6936_o ? n7227_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7305_o = n6936_o ? n7228_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7306_o = n6936_o ? n7230_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7308_o = n6936_o ? n7232_o : 2'b00;
  /* TG68KdotC_Kernel.vhd:3008:33  */
  assign n7309_o = n6936_o ? n7233_o : n7256_o;
  /* TG68KdotC_Kernel.vhd:3007:25  */
  assign n7311_o = n2185_o == 4'b1110;
  /* TG68KdotC_Kernel.vhd:3117:39  */
  assign n7312_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:3117:57  */
  assign n7313_o = opcode[8:6];
  /* TG68KdotC_Kernel.vhd:3117:69  */
  assign n7315_o = n7313_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:3117:47  */
  assign n7316_o = n7315_o & n7312_o;
  /* TG68KdotC_Kernel.vhd:3118:50  */
  assign n7317_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:3118:62  */
  assign n7319_o = n7317_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:3118:79  */
  assign n7320_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:3118:91  */
  assign n7322_o = n7320_o != 3'b011;
  /* TG68KdotC_Kernel.vhd:3118:69  */
  assign n7323_o = n7322_o & n7319_o;
  /* TG68KdotC_Kernel.vhd:3119:51  */
  assign n7324_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:3119:63  */
  assign n7326_o = n7324_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:3119:80  */
  assign n7327_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:3119:92  */
  assign n7329_o = n7327_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:3119:71  */
  assign n7330_o = n7326_o | n7329_o;
  /* TG68KdotC_Kernel.vhd:3118:99  */
  assign n7331_o = n7330_o & n7323_o;
  /* TG68KdotC_Kernel.vhd:3120:58  */
  assign n7332_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:3120:71  */
  assign n7334_o = n7332_o != 3'b000;
  /* TG68KdotC_Kernel.vhd:3122:74  */
  assign n7335_o = opcode[5];
  /* TG68KdotC_Kernel.vhd:3122:77  */
  assign n7336_o = ~n7335_o;
  /* TG68KdotC_Kernel.vhd:3122:92  */
  assign n7337_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:3122:104  */
  assign n7339_o = n7337_o != 2'b01;
  /* TG68KdotC_Kernel.vhd:3122:82  */
  assign n7340_o = n7339_o & n7336_o;
  /* TG68KdotC_Kernel.vhd:3122:65  */
  assign n7343_o = n7340_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3122:65  */
  assign n7346_o = n7340_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3121:57  */
  assign n7348_o = svmode ? n7343_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3121:57  */
  assign n7351_o = svmode ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3121:57  */
  assign n7353_o = svmode ? n7346_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3136:57  */
  assign n7356_o = svmode ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3136:57  */
  assign n7359_o = svmode ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3120:49  */
  assign n7361_o = n7334_o ? n7348_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3120:49  */
  assign n7362_o = n7334_o ? n7351_o : n7356_o;
  /* TG68KdotC_Kernel.vhd:3120:49  */
  assign n7363_o = n7334_o ? n7353_o : n7359_o;
  /* TG68KdotC_Kernel.vhd:3118:41  */
  assign n7365_o = n7331_o ? n7361_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3118:41  */
  assign n7367_o = n7331_o ? n7362_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3118:41  */
  assign n7369_o = n7331_o ? n7363_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3148:42  */
  assign n7370_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:3148:60  */
  assign n7371_o = opcode[8:6];
  /* TG68KdotC_Kernel.vhd:3148:72  */
  assign n7373_o = n7371_o == 3'b101;
  /* TG68KdotC_Kernel.vhd:3148:50  */
  assign n7374_o = n7373_o & n7370_o;
  /* TG68KdotC_Kernel.vhd:3149:50  */
  assign n7375_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:3149:62  */
  assign n7377_o = n7375_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:3149:79  */
  assign n7378_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:3149:91  */
  assign n7380_o = n7378_o != 3'b100;
  /* TG68KdotC_Kernel.vhd:3149:69  */
  assign n7381_o = n7380_o & n7377_o;
  /* TG68KdotC_Kernel.vhd:3150:51  */
  assign n7382_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:3150:63  */
  assign n7384_o = n7382_o != 3'b111;
  /* TG68KdotC_Kernel.vhd:3150:81  */
  assign n7385_o = opcode[2:1];
  /* TG68KdotC_Kernel.vhd:3150:93  */
  assign n7387_o = n7385_o != 2'b11;
  /* TG68KdotC_Kernel.vhd:3151:50  */
  assign n7388_o = opcode[2:0];
  /* TG68KdotC_Kernel.vhd:3151:62  */
  assign n7390_o = n7388_o != 3'b101;
  /* TG68KdotC_Kernel.vhd:3150:100  */
  assign n7391_o = n7390_o & n7387_o;
  /* TG68KdotC_Kernel.vhd:3150:71  */
  assign n7392_o = n7384_o | n7391_o;
  /* TG68KdotC_Kernel.vhd:3149:99  */
  assign n7393_o = n7392_o & n7381_o;
  /* TG68KdotC_Kernel.vhd:3152:58  */
  assign n7394_o = opcode[5:1];
  /* TG68KdotC_Kernel.vhd:3152:70  */
  assign n7396_o = n7394_o != 5'b11110;
  /* TG68KdotC_Kernel.vhd:3153:66  */
  assign n7397_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:3153:79  */
  assign n7399_o = n7397_o == 3'b001;
  /* TG68KdotC_Kernel.vhd:3153:95  */
  assign n7400_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:3153:108  */
  assign n7402_o = n7400_o == 3'b010;
  /* TG68KdotC_Kernel.vhd:3153:86  */
  assign n7403_o = n7399_o | n7402_o;
  /* TG68KdotC_Kernel.vhd:3155:82  */
  assign n7404_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:3155:94  */
  assign n7406_o = n7404_o == 3'b101;
  /* TG68KdotC_Kernel.vhd:3155:73  */
  assign n7409_o = n7406_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3155:73  */
  assign n7412_o = n7406_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3154:65  */
  assign n7414_o = svmode ? n7409_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3154:65  */
  assign n7417_o = svmode ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3154:65  */
  assign n7419_o = svmode ? n7412_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3168:65  */
  assign n7422_o = svmode ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3168:65  */
  assign n7425_o = svmode ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3153:57  */
  assign n7427_o = n7403_o ? n7414_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3153:57  */
  assign n7428_o = n7403_o ? n7417_o : n7422_o;
  /* TG68KdotC_Kernel.vhd:3153:57  */
  assign n7429_o = n7403_o ? n7419_o : n7425_o;
  /* TG68KdotC_Kernel.vhd:3152:49  */
  assign n7431_o = n7396_o ? n7427_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3152:49  */
  assign n7433_o = n7396_o ? n7428_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3152:49  */
  assign n7435_o = n7396_o ? n7429_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3149:41  */
  assign n7437_o = n7393_o ? n7431_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3149:41  */
  assign n7439_o = n7393_o ? n7433_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3149:41  */
  assign n7441_o = n7393_o ? n7435_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3148:33  */
  assign n7443_o = n7374_o ? n7437_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3148:33  */
  assign n7445_o = n7374_o ? n7439_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3148:33  */
  assign n7447_o = n7374_o ? n7441_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3117:33  */
  assign n7448_o = n7316_o ? n7365_o : n7443_o;
  /* TG68KdotC_Kernel.vhd:3117:33  */
  assign n7449_o = n7316_o ? n7367_o : n7445_o;
  /* TG68KdotC_Kernel.vhd:3117:33  */
  assign n7450_o = n7316_o ? n7369_o : n7447_o;
  /* TG68KdotC_Kernel.vhd:3116:25  */
  assign n7452_o = n2185_o == 4'b1111;
  assign n7453_o = {n7452_o, n7311_o, n6933_o, n6672_o, n6459_o, n6457_o, n6340_o, n6017_o, n5994_o, n5932_o, n5712_o, n3355_o, n3141_o};
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7454_o = make_berr;
      13'b0100000000000: n7454_o = make_berr;
      13'b0010000000000: n7454_o = make_berr;
      13'b0001000000000: n7454_o = make_berr;
      13'b0000100000000: n7454_o = make_berr;
      13'b0000010000000: n7454_o = make_berr;
      13'b0000001000000: n7454_o = make_berr;
      13'b0000000100000: n7454_o = make_berr;
      13'b0000000010000: n7454_o = make_berr;
      13'b0000000001000: n7454_o = n5905_o;
      13'b0000000000100: n7454_o = n5603_o;
      13'b0000000000010: n7454_o = make_berr;
      13'b0000000000001: n7454_o = make_berr;
      default: n7454_o = make_berr;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7456_o = n1921_o;
      13'b0100000000000: n7456_o = n6954_o;
      13'b0010000000000: n7456_o = n6896_o;
      13'b0001000000000: n7456_o = n6474_o;
      13'b0000100000000: n7456_o = n1921_o;
      13'b0000010000000: n7456_o = n6381_o;
      13'b0000001000000: n7456_o = n6301_o;
      13'b0000000100000: n7456_o = n6001_o;
      13'b0000000010000: n7456_o = 2'b10;
      13'b0000000001000: n7456_o = n5906_o;
      13'b0000000000100: n7456_o = n5604_o;
      13'b0000000000010: n7456_o = n3314_o;
      13'b0000000000001: n7456_o = n3080_o;
      default: n7456_o = n1921_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7457_o = datatype;
      13'b0100000000000: n7457_o = datatype;
      13'b0010000000000: n7457_o = datatype;
      13'b0001000000000: n7457_o = datatype;
      13'b0000100000000: n7457_o = datatype;
      13'b0000010000000: n7457_o = datatype;
      13'b0000001000000: n7457_o = n6302_o;
      13'b0000000100000: n7457_o = datatype;
      13'b0000000010000: n7457_o = datatype;
      13'b0000000001000: n7457_o = datatype;
      13'b0000000000100: n7457_o = datatype;
      13'b0000000000010: n7457_o = datatype;
      13'b0000000000001: n7457_o = datatype;
      default: n7457_o = datatype;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7458_o = n2026_o;
      13'b0100000000000: n7458_o = n7266_o;
      13'b0010000000000: n7458_o = n6897_o;
      13'b0001000000000: n7458_o = n6639_o;
      13'b0000100000000: n7458_o = n2026_o;
      13'b0000010000000: n7458_o = n2026_o;
      13'b0000001000000: n7458_o = n6049_o;
      13'b0000000100000: n7458_o = n2026_o;
      13'b0000000010000: n7458_o = n5983_o;
      13'b0000000001000: n7458_o = n5907_o;
      13'b0000000000100: n7458_o = n5605_o;
      13'b0000000000010: n7458_o = n3304_o;
      13'b0000000000001: n7458_o = n3081_o;
      default: n7458_o = n2026_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7459_o = n2148_o;
      13'b0100000000000: n7459_o = n2148_o;
      13'b0010000000000: n7459_o = n2148_o;
      13'b0001000000000: n7459_o = n2148_o;
      13'b0000100000000: n7459_o = n2148_o;
      13'b0000010000000: n7459_o = n2148_o;
      13'b0000001000000: n7459_o = n2148_o;
      13'b0000000100000: n7459_o = n2148_o;
      13'b0000000010000: n7459_o = n2148_o;
      13'b0000000001000: n7459_o = n2148_o;
      13'b0000000000100: n7459_o = n5606_o;
      13'b0000000000010: n7459_o = n2148_o;
      13'b0000000000001: n7459_o = n2148_o;
      default: n7459_o = n2148_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7461_o = 1'b0;
      13'b0100000000000: n7461_o = 1'b0;
      13'b0010000000000: n7461_o = n6899_o;
      13'b0001000000000: n7461_o = 1'b0;
      13'b0000100000000: n7461_o = 1'b0;
      13'b0000010000000: n7461_o = 1'b0;
      13'b0000001000000: n7461_o = n6305_o;
      13'b0000000100000: n7461_o = 1'b0;
      13'b0000000010000: n7461_o = 1'b0;
      13'b0000000001000: n7461_o = 1'b0;
      13'b0000000000100: n7461_o = 1'b0;
      13'b0000000000010: n7461_o = 1'b0;
      13'b0000000000001: n7461_o = 1'b0;
      default: n7461_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7462_o = n2151_o;
      13'b0100000000000: n7462_o = n2151_o;
      13'b0010000000000: n7462_o = n2151_o;
      13'b0001000000000: n7462_o = n2151_o;
      13'b0000100000000: n7462_o = n2151_o;
      13'b0000010000000: n7462_o = n2151_o;
      13'b0000001000000: n7462_o = n2151_o;
      13'b0000000100000: n7462_o = n2151_o;
      13'b0000000010000: n7462_o = n2151_o;
      13'b0000000001000: n7462_o = n2151_o;
      13'b0000000000100: n7462_o = n5607_o;
      13'b0000000000010: n7462_o = n3305_o;
      13'b0000000000001: n7462_o = n2151_o;
      default: n7462_o = n2151_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7464_o = 1'b0;
      13'b0100000000000: n7464_o = n7269_o;
      13'b0010000000000: n7464_o = 1'b0;
      13'b0001000000000: n7464_o = 1'b0;
      13'b0000100000000: n7464_o = 1'b0;
      13'b0000010000000: n7464_o = 1'b0;
      13'b0000001000000: n7464_o = 1'b0;
      13'b0000000100000: n7464_o = 1'b0;
      13'b0000000010000: n7464_o = 1'b0;
      13'b0000000001000: n7464_o = n5909_o;
      13'b0000000000100: n7464_o = 1'b0;
      13'b0000000000010: n7464_o = 1'b0;
      13'b0000000000001: n7464_o = 1'b0;
      default: n7464_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7466_o = 1'b0;
      13'b0100000000000: n7466_o = n7271_o;
      13'b0010000000000: n7466_o = 1'b0;
      13'b0001000000000: n7466_o = 1'b0;
      13'b0000100000000: n7466_o = 1'b0;
      13'b0000010000000: n7466_o = 1'b0;
      13'b0000001000000: n7466_o = n6307_o;
      13'b0000000100000: n7466_o = 1'b0;
      13'b0000000010000: n7466_o = 1'b0;
      13'b0000000001000: n7466_o = n5910_o;
      13'b0000000000100: n7466_o = n5609_o;
      13'b0000000000010: n7466_o = 1'b0;
      13'b0000000000001: n7466_o = n3083_o;
      default: n7466_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7467_o = n2015_o;
      13'b0100000000000: n7467_o = n2015_o;
      13'b0010000000000: n7467_o = n2015_o;
      13'b0001000000000: n7467_o = n2015_o;
      13'b0000100000000: n7467_o = n2015_o;
      13'b0000010000000: n7467_o = n2015_o;
      13'b0000001000000: n7467_o = n2015_o;
      13'b0000000100000: n7467_o = n2015_o;
      13'b0000000010000: n7467_o = n5973_o;
      13'b0000000001000: n7467_o = n2015_o;
      13'b0000000000100: n7467_o = n5610_o;
      13'b0000000000010: n7467_o = n2015_o;
      13'b0000000000001: n7467_o = n2015_o;
      default: n7467_o = n2015_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7469_o = 1'b0;
      13'b0100000000000: n7469_o = 1'b0;
      13'b0010000000000: n7469_o = 1'b0;
      13'b0001000000000: n7469_o = 1'b0;
      13'b0000100000000: n7469_o = 1'b0;
      13'b0000010000000: n7469_o = 1'b0;
      13'b0000001000000: n7469_o = 1'b0;
      13'b0000000100000: n7469_o = 1'b0;
      13'b0000000010000: n7469_o = n5986_o;
      13'b0000000001000: n7469_o = 1'b0;
      13'b0000000000100: n7469_o = n5612_o;
      13'b0000000000010: n7469_o = 1'b0;
      13'b0000000000001: n7469_o = 1'b0;
      default: n7469_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7471_o = 1'b0;
      13'b0100000000000: n7471_o = 1'b0;
      13'b0010000000000: n7471_o = 1'b0;
      13'b0001000000000: n7471_o = 1'b0;
      13'b0000100000000: n7471_o = 1'b0;
      13'b0000010000000: n7471_o = 1'b0;
      13'b0000001000000: n7471_o = 1'b0;
      13'b0000000100000: n7471_o = 1'b0;
      13'b0000000010000: n7471_o = 1'b0;
      13'b0000000001000: n7471_o = 1'b0;
      13'b0000000000100: n7471_o = n5614_o;
      13'b0000000000010: n7471_o = 1'b0;
      13'b0000000000001: n7471_o = 1'b0;
      default: n7471_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7473_o = 1'b0;
      13'b0100000000000: n7473_o = n7273_o;
      13'b0010000000000: n7473_o = 1'b0;
      13'b0001000000000: n7473_o = 1'b0;
      13'b0000100000000: n7473_o = 1'b0;
      13'b0000010000000: n7473_o = 1'b0;
      13'b0000001000000: n7473_o = 1'b0;
      13'b0000000100000: n7473_o = 1'b0;
      13'b0000000010000: n7473_o = 1'b0;
      13'b0000000001000: n7473_o = 1'b0;
      13'b0000000000100: n7473_o = n5615_o;
      13'b0000000000010: n7473_o = 1'b0;
      13'b0000000000001: n7473_o = 1'b0;
      default: n7473_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7475_o = 1'b0;
      13'b0100000000000: n7475_o = 1'b0;
      13'b0010000000000: n7475_o = n6901_o;
      13'b0001000000000: n7475_o = n6641_o;
      13'b0000100000000: n7475_o = 1'b0;
      13'b0000010000000: n7475_o = n6425_o;
      13'b0000001000000: n7475_o = 1'b0;
      13'b0000000100000: n7475_o = 1'b0;
      13'b0000000010000: n7475_o = 1'b0;
      13'b0000000001000: n7475_o = 1'b0;
      13'b0000000000100: n7475_o = n5616_o;
      13'b0000000000010: n7475_o = n3318_o;
      13'b0000000000001: n7475_o = 1'b0;
      default: n7475_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7477_o = 1'b0;
      13'b0100000000000: n7477_o = n7275_o;
      13'b0010000000000: n7477_o = n6903_o;
      13'b0001000000000: n7477_o = n6643_o;
      13'b0000100000000: n7477_o = 1'b0;
      13'b0000010000000: n7477_o = n6427_o;
      13'b0000001000000: n7477_o = n6308_o;
      13'b0000000100000: n7477_o = 1'b0;
      13'b0000000010000: n7477_o = 1'b0;
      13'b0000000001000: n7477_o = 1'b0;
      13'b0000000000100: n7477_o = n5617_o;
      13'b0000000000010: n7477_o = n3321_o;
      13'b0000000000001: n7477_o = 1'b0;
      default: n7477_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7479_o = 1'b0;
      13'b0100000000000: n7479_o = n7277_o;
      13'b0010000000000: n7479_o = 1'b0;
      13'b0001000000000: n7479_o = 1'b0;
      13'b0000100000000: n7479_o = 1'b0;
      13'b0000010000000: n7479_o = 1'b0;
      13'b0000001000000: n7479_o = 1'b0;
      13'b0000000100000: n7479_o = 1'b0;
      13'b0000000010000: n7479_o = 1'b0;
      13'b0000000001000: n7479_o = 1'b0;
      13'b0000000000100: n7479_o = 1'b0;
      13'b0000000000010: n7479_o = 1'b0;
      13'b0000000000001: n7479_o = 1'b0;
      default: n7479_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7481_o = 1'b0;
      13'b0100000000000: n7481_o = n7279_o;
      13'b0010000000000: n7481_o = 1'b0;
      13'b0001000000000: n7481_o = 1'b0;
      13'b0000100000000: n7481_o = 1'b0;
      13'b0000010000000: n7481_o = 1'b0;
      13'b0000001000000: n7481_o = 1'b0;
      13'b0000000100000: n7481_o = 1'b0;
      13'b0000000010000: n7481_o = 1'b0;
      13'b0000000001000: n7481_o = 1'b0;
      13'b0000000000100: n7481_o = n5619_o;
      13'b0000000000010: n7481_o = 1'b0;
      13'b0000000000001: n7481_o = n3085_o;
      default: n7481_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7483_o = 1'b0;
      13'b0100000000000: n7483_o = 1'b0;
      13'b0010000000000: n7483_o = n6905_o;
      13'b0001000000000: n7483_o = n6645_o;
      13'b0000100000000: n7483_o = 1'b0;
      13'b0000010000000: n7483_o = n6429_o;
      13'b0000001000000: n7483_o = 1'b0;
      13'b0000000100000: n7483_o = 1'b0;
      13'b0000000010000: n7483_o = 1'b0;
      13'b0000000001000: n7483_o = 1'b0;
      13'b0000000000100: n7483_o = n5621_o;
      13'b0000000000010: n7483_o = n3323_o;
      13'b0000000000001: n7483_o = 1'b0;
      default: n7483_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7485_o = 1'b0;
      13'b0100000000000: n7485_o = n7281_o;
      13'b0010000000000: n7485_o = 1'b0;
      13'b0001000000000: n7485_o = 1'b0;
      13'b0000100000000: n7485_o = 1'b0;
      13'b0000010000000: n7485_o = 1'b0;
      13'b0000001000000: n7485_o = 1'b0;
      13'b0000000100000: n7485_o = 1'b0;
      13'b0000000010000: n7485_o = 1'b0;
      13'b0000000001000: n7485_o = 1'b0;
      13'b0000000000100: n7485_o = n5623_o;
      13'b0000000000010: n7485_o = 1'b0;
      13'b0000000000001: n7485_o = 1'b0;
      default: n7485_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7487_o = 1'b0;
      13'b0100000000000: n7487_o = 1'b0;
      13'b0010000000000: n7487_o = n6906_o;
      13'b0001000000000: n7487_o = n6647_o;
      13'b0000100000000: n7487_o = 1'b0;
      13'b0000010000000: n7487_o = n6431_o;
      13'b0000001000000: n7487_o = n6309_o;
      13'b0000000100000: n7487_o = n6004_o;
      13'b0000000010000: n7487_o = 1'b0;
      13'b0000000001000: n7487_o = 1'b0;
      13'b0000000000100: n7487_o = n5624_o;
      13'b0000000000010: n7487_o = n3325_o;
      13'b0000000000001: n7487_o = n3087_o;
      default: n7487_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7488_o = n1900_o;
      13'b0100000000000: n7488_o = n6958_o;
      13'b0010000000000: n7488_o = n1900_o;
      13'b0001000000000: n7488_o = n1900_o;
      13'b0000100000000: n7488_o = n1900_o;
      13'b0000010000000: n7488_o = n1900_o;
      13'b0000001000000: n7488_o = n1900_o;
      13'b0000000100000: n7488_o = n1900_o;
      13'b0000000010000: n7488_o = n1900_o;
      13'b0000000001000: n7488_o = n1900_o;
      13'b0000000000100: n7488_o = n1900_o;
      13'b0000000000010: n7488_o = n1900_o;
      13'b0000000000001: n7488_o = n1900_o;
      default: n7488_o = n1900_o;
    endcase
  assign n7489_o = n5625_o[3:0];
  assign n7490_o = n1904_o[3:0];
  assign n7491_o = n1905_o[3:0];
  /* TG68KdotC_Kernel.vhd:1495:17  */
  assign n7492_o = n1902_o ? n7490_o : n7491_o;
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7493_o = n7492_o;
      13'b0100000000000: n7493_o = n7286_o;
      13'b0010000000000: n7493_o = n7492_o;
      13'b0001000000000: n7493_o = n7492_o;
      13'b0000100000000: n7493_o = n7492_o;
      13'b0000010000000: n7493_o = n7492_o;
      13'b0000001000000: n7493_o = n7492_o;
      13'b0000000100000: n7493_o = n7492_o;
      13'b0000000010000: n7493_o = n7492_o;
      13'b0000000001000: n7493_o = n7492_o;
      13'b0000000000100: n7493_o = n7489_o;
      13'b0000000000010: n7493_o = n7492_o;
      13'b0000000000001: n7493_o = n7492_o;
      default: n7493_o = n7492_o;
    endcase
  assign n7494_o = n5625_o[5:4];
  assign n7495_o = n1904_o[5:4];
  assign n7496_o = n1905_o[5:4];
  /* TG68KdotC_Kernel.vhd:1495:17  */
  assign n7497_o = n1902_o ? n7495_o : n7496_o;
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7498_o = n7497_o;
      13'b0100000000000: n7498_o = n7497_o;
      13'b0010000000000: n7498_o = n7497_o;
      13'b0001000000000: n7498_o = n7497_o;
      13'b0000100000000: n7498_o = n7497_o;
      13'b0000010000000: n7498_o = n7497_o;
      13'b0000001000000: n7498_o = n7497_o;
      13'b0000000100000: n7498_o = n7497_o;
      13'b0000000010000: n7498_o = n7497_o;
      13'b0000000001000: n7498_o = n7497_o;
      13'b0000000000100: n7498_o = n7494_o;
      13'b0000000000010: n7498_o = n7497_o;
      13'b0000000000001: n7498_o = n7497_o;
      default: n7498_o = n7497_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7500_o = 1'b0;
      13'b0100000000000: n7500_o = 1'b0;
      13'b0010000000000: n7500_o = 1'b0;
      13'b0001000000000: n7500_o = 1'b0;
      13'b0000100000000: n7500_o = 1'b0;
      13'b0000010000000: n7500_o = 1'b0;
      13'b0000001000000: n7500_o = 1'b0;
      13'b0000000100000: n7500_o = 1'b0;
      13'b0000000010000: n7500_o = 1'b0;
      13'b0000000001000: n7500_o = 1'b0;
      13'b0000000000100: n7500_o = n5627_o;
      13'b0000000000010: n7500_o = 1'b0;
      13'b0000000000001: n7500_o = 1'b0;
      default: n7500_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7501_o = n2154_o;
      13'b0100000000000: n7501_o = n2154_o;
      13'b0010000000000: n7501_o = n2154_o;
      13'b0001000000000: n7501_o = n2154_o;
      13'b0000100000000: n7501_o = n2154_o;
      13'b0000010000000: n7501_o = n2154_o;
      13'b0000001000000: n7501_o = n6310_o;
      13'b0000000100000: n7501_o = n2154_o;
      13'b0000000010000: n7501_o = n2154_o;
      13'b0000000001000: n7501_o = n2154_o;
      13'b0000000000100: n7501_o = n5628_o;
      13'b0000000000010: n7501_o = n2154_o;
      13'b0000000000001: n7501_o = n3088_o;
      default: n7501_o = n2154_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7504_o = n7448_o;
      13'b0100000000000: n7504_o = n7288_o;
      13'b0010000000000: n7504_o = n6907_o;
      13'b0001000000000: n7504_o = n6648_o;
      13'b0000100000000: n7504_o = 1'b0;
      13'b0000010000000: n7504_o = n6434_o;
      13'b0000001000000: n7504_o = n6311_o;
      13'b0000000100000: n7504_o = n6007_o;
      13'b0000000010000: n7504_o = 1'b0;
      13'b0000000001000: n7504_o = n5911_o;
      13'b0000000000100: n7504_o = n5629_o;
      13'b0000000000010: n7504_o = n3328_o;
      13'b0000000000001: n7504_o = n3090_o;
      default: n7504_o = 1'b1;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7506_o = n7449_o;
      13'b0100000000000: n7506_o = 1'b0;
      13'b0010000000000: n7506_o = 1'b0;
      13'b0001000000000: n7506_o = 1'b0;
      13'b0000100000000: n7506_o = 1'b0;
      13'b0000010000000: n7506_o = 1'b0;
      13'b0000001000000: n7506_o = 1'b0;
      13'b0000000100000: n7506_o = 1'b0;
      13'b0000000010000: n7506_o = 1'b0;
      13'b0000000001000: n7506_o = 1'b0;
      13'b0000000000100: n7506_o = n5631_o;
      13'b0000000000010: n7506_o = 1'b0;
      13'b0000000000001: n7506_o = n3092_o;
      default: n7506_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7509_o = 1'b0;
      13'b0100000000000: n7509_o = 1'b0;
      13'b0010000000000: n7509_o = 1'b0;
      13'b0001000000000: n7509_o = 1'b0;
      13'b0000100000000: n7509_o = 1'b1;
      13'b0000010000000: n7509_o = 1'b0;
      13'b0000001000000: n7509_o = 1'b0;
      13'b0000000100000: n7509_o = 1'b0;
      13'b0000000010000: n7509_o = 1'b0;
      13'b0000000001000: n7509_o = 1'b0;
      13'b0000000000100: n7509_o = 1'b0;
      13'b0000000000010: n7509_o = 1'b0;
      13'b0000000000001: n7509_o = 1'b0;
      default: n7509_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7511_o = n7450_o;
      13'b0100000000000: n7511_o = 1'b0;
      13'b0010000000000: n7511_o = 1'b0;
      13'b0001000000000: n7511_o = 1'b0;
      13'b0000100000000: n7511_o = 1'b0;
      13'b0000010000000: n7511_o = 1'b0;
      13'b0000001000000: n7511_o = 1'b0;
      13'b0000000100000: n7511_o = 1'b0;
      13'b0000000010000: n7511_o = 1'b0;
      13'b0000000001000: n7511_o = 1'b0;
      13'b0000000000100: n7511_o = 1'b0;
      13'b0000000000010: n7511_o = 1'b0;
      13'b0000000000001: n7511_o = 1'b0;
      default: n7511_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7513_o = 1'b0;
      13'b0100000000000: n7513_o = 1'b0;
      13'b0010000000000: n7513_o = 1'b0;
      13'b0001000000000: n7513_o = 1'b0;
      13'b0000100000000: n7513_o = 1'b0;
      13'b0000010000000: n7513_o = 1'b0;
      13'b0000001000000: n7513_o = 1'b0;
      13'b0000000100000: n7513_o = 1'b0;
      13'b0000000010000: n7513_o = 1'b0;
      13'b0000000001000: n7513_o = 1'b0;
      13'b0000000000100: n7513_o = n5633_o;
      13'b0000000000010: n7513_o = 1'b0;
      13'b0000000000001: n7513_o = 1'b0;
      default: n7513_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7515_o = 1'b0;
      13'b0100000000000: n7515_o = 1'b0;
      13'b0010000000000: n7515_o = 1'b0;
      13'b0001000000000: n7515_o = 1'b0;
      13'b0000100000000: n7515_o = 1'b0;
      13'b0000010000000: n7515_o = 1'b0;
      13'b0000001000000: n7515_o = 1'b0;
      13'b0000000100000: n7515_o = 1'b0;
      13'b0000000010000: n7515_o = 1'b0;
      13'b0000000001000: n7515_o = n5913_o;
      13'b0000000000100: n7515_o = n5635_o;
      13'b0000000000010: n7515_o = 1'b0;
      13'b0000000000001: n7515_o = 1'b0;
      default: n7515_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7520_o = 1'b1;
      13'b0100000000000: n7520_o = n7290_o;
      13'b0010000000000: n7520_o = n6908_o;
      13'b0001000000000: n7520_o = n6649_o;
      13'b0000100000000: n7520_o = 1'b1;
      13'b0000010000000: n7520_o = n6437_o;
      13'b0000001000000: n7520_o = n6312_o;
      13'b0000000100000: n7520_o = n6010_o;
      13'b0000000010000: n7520_o = 1'b0;
      13'b0000000001000: n7520_o = n5914_o;
      13'b0000000000100: n7520_o = n5636_o;
      13'b0000000000010: n7520_o = n3331_o;
      13'b0000000000001: n7520_o = n3094_o;
      default: n7520_o = 1'b1;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7522_o = 1'b0;
      13'b0100000000000: n7522_o = 1'b0;
      13'b0010000000000: n7522_o = 1'b0;
      13'b0001000000000: n7522_o = 1'b0;
      13'b0000100000000: n7522_o = 1'b0;
      13'b0000010000000: n7522_o = 1'b0;
      13'b0000001000000: n7522_o = 1'b0;
      13'b0000000100000: n7522_o = 1'b0;
      13'b0000000010000: n7522_o = 1'b0;
      13'b0000000001000: n7522_o = 1'b0;
      13'b0000000000100: n7522_o = n5638_o;
      13'b0000000000010: n7522_o = 1'b0;
      13'b0000000000001: n7522_o = 1'b0;
      default: n7522_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7524_o = 1'b0;
      13'b0100000000000: n7524_o = n7292_o;
      13'b0010000000000: n7524_o = n6910_o;
      13'b0001000000000: n7524_o = n6650_o;
      13'b0000100000000: n7524_o = 1'b0;
      13'b0000010000000: n7524_o = n6440_o;
      13'b0000001000000: n7524_o = n6314_o;
      13'b0000000100000: n7524_o = 1'b0;
      13'b0000000010000: n7524_o = 1'b0;
      13'b0000000001000: n7524_o = n5915_o;
      13'b0000000000100: n7524_o = n5639_o;
      13'b0000000000010: n7524_o = n3334_o;
      13'b0000000000001: n7524_o = n3096_o;
      default: n7524_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7526_o = 1'b0;
      13'b0100000000000: n7526_o = 1'b0;
      13'b0010000000000: n7526_o = n6912_o;
      13'b0001000000000: n7526_o = n6652_o;
      13'b0000100000000: n7526_o = 1'b0;
      13'b0000010000000: n7526_o = n6442_o;
      13'b0000001000000: n7526_o = n6316_o;
      13'b0000000100000: n7526_o = 1'b0;
      13'b0000000010000: n7526_o = 1'b0;
      13'b0000000001000: n7526_o = 1'b0;
      13'b0000000000100: n7526_o = 1'b0;
      13'b0000000000010: n7526_o = 1'b0;
      13'b0000000000001: n7526_o = 1'b0;
      default: n7526_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7528_o = 1'b0;
      13'b0100000000000: n7528_o = 1'b0;
      13'b0010000000000: n7528_o = n6914_o;
      13'b0001000000000: n7528_o = 1'b0;
      13'b0000100000000: n7528_o = 1'b0;
      13'b0000010000000: n7528_o = n6444_o;
      13'b0000001000000: n7528_o = n6318_o;
      13'b0000000100000: n7528_o = 1'b0;
      13'b0000000010000: n7528_o = 1'b0;
      13'b0000000001000: n7528_o = 1'b0;
      13'b0000000000100: n7528_o = 1'b0;
      13'b0000000000010: n7528_o = 1'b0;
      13'b0000000000001: n7528_o = 1'b0;
      default: n7528_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7530_o = 1'b0;
      13'b0100000000000: n7530_o = 1'b0;
      13'b0010000000000: n7530_o = 1'b0;
      13'b0001000000000: n7530_o = 1'b0;
      13'b0000100000000: n7530_o = 1'b0;
      13'b0000010000000: n7530_o = 1'b0;
      13'b0000001000000: n7530_o = 1'b0;
      13'b0000000100000: n7530_o = 1'b0;
      13'b0000000010000: n7530_o = 1'b0;
      13'b0000000001000: n7530_o = 1'b0;
      13'b0000000000100: n7530_o = 1'b0;
      13'b0000000000010: n7530_o = 1'b0;
      13'b0000000000001: n7530_o = n3098_o;
      default: n7530_o = 1'b0;
    endcase
  assign n7531_o = n1909_o[0];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7532_o = n7531_o;
      13'b0100000000000: n7532_o = n7531_o;
      13'b0010000000000: n7532_o = n7531_o;
      13'b0001000000000: n7532_o = n7531_o;
      13'b0000100000000: n7532_o = n7531_o;
      13'b0000010000000: n7532_o = n7531_o;
      13'b0000001000000: n7532_o = n7531_o;
      13'b0000000100000: n7532_o = n7531_o;
      13'b0000000010000: n7532_o = n7531_o;
      13'b0000000001000: n7532_o = n7531_o;
      13'b0000000000100: n7532_o = n5645_o;
      13'b0000000000010: n7532_o = n7531_o;
      13'b0000000000001: n7532_o = n7531_o;
      default: n7532_o = n7531_o;
    endcase
  assign n7533_o = n1909_o[19:17];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7534_o = n7533_o;
      13'b0100000000000: n7534_o = n7533_o;
      13'b0010000000000: n7534_o = n7533_o;
      13'b0001000000000: n7534_o = n7533_o;
      13'b0000100000000: n7534_o = n7533_o;
      13'b0000010000000: n7534_o = n7533_o;
      13'b0000001000000: n7534_o = n7533_o;
      13'b0000000100000: n7534_o = n7533_o;
      13'b0000000010000: n7534_o = n7533_o;
      13'b0000000001000: n7534_o = n7533_o;
      13'b0000000000100: n7534_o = n7533_o;
      13'b0000000000010: n7534_o = n7533_o;
      13'b0000000000001: n7534_o = n3102_o;
      default: n7534_o = n7533_o;
    endcase
  assign n7535_o = n1909_o[24];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7536_o = n7535_o;
      13'b0100000000000: n7536_o = n7294_o;
      13'b0010000000000: n7536_o = n6707_o;
      13'b0001000000000: n7536_o = n7535_o;
      13'b0000100000000: n7536_o = n7535_o;
      13'b0000010000000: n7536_o = n7535_o;
      13'b0000001000000: n7536_o = n7535_o;
      13'b0000000100000: n7536_o = n7535_o;
      13'b0000000010000: n7536_o = n7535_o;
      13'b0000000001000: n7536_o = n7535_o;
      13'b0000000000100: n7536_o = n5647_o;
      13'b0000000000010: n7536_o = n7535_o;
      13'b0000000000001: n7536_o = n7535_o;
      default: n7536_o = n7535_o;
    endcase
  assign n7537_o = n1909_o[26];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7538_o = n7537_o;
      13'b0100000000000: n7538_o = n7537_o;
      13'b0010000000000: n7538_o = n7537_o;
      13'b0001000000000: n7538_o = n7537_o;
      13'b0000100000000: n7538_o = n7537_o;
      13'b0000010000000: n7538_o = n7537_o;
      13'b0000001000000: n7538_o = n7537_o;
      13'b0000000100000: n7538_o = n7537_o;
      13'b0000000010000: n7538_o = n7537_o;
      13'b0000000001000: n7538_o = n7537_o;
      13'b0000000000100: n7538_o = n7537_o;
      13'b0000000000010: n7538_o = n7537_o;
      13'b0000000000001: n7538_o = n3104_o;
      default: n7538_o = n7537_o;
    endcase
  assign n7539_o = n1909_o[29];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7540_o = n7539_o;
      13'b0100000000000: n7540_o = n7296_o;
      13'b0010000000000: n7540_o = n7539_o;
      13'b0001000000000: n7540_o = n7539_o;
      13'b0000100000000: n7540_o = n7539_o;
      13'b0000010000000: n7540_o = n7539_o;
      13'b0000001000000: n7540_o = n7539_o;
      13'b0000000100000: n7540_o = n7539_o;
      13'b0000000010000: n7540_o = n7539_o;
      13'b0000000001000: n7540_o = n7539_o;
      13'b0000000000100: n7540_o = n7539_o;
      13'b0000000000010: n7540_o = n7539_o;
      13'b0000000000001: n7540_o = n7539_o;
      default: n7540_o = n7539_o;
    endcase
  assign n7541_o = n1909_o[34];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7542_o = n7541_o;
      13'b0100000000000: n7542_o = n7541_o;
      13'b0010000000000: n7542_o = n6918_o;
      13'b0001000000000: n7542_o = n7541_o;
      13'b0000100000000: n7542_o = n7541_o;
      13'b0000010000000: n7542_o = n7541_o;
      13'b0000001000000: n7542_o = n7541_o;
      13'b0000000100000: n7542_o = n7541_o;
      13'b0000000010000: n7542_o = n7541_o;
      13'b0000000001000: n7542_o = n7541_o;
      13'b0000000000100: n7542_o = n5649_o;
      13'b0000000000010: n7542_o = n7541_o;
      13'b0000000000001: n7542_o = n7541_o;
      default: n7542_o = n7541_o;
    endcase
  assign n7543_o = n1909_o[36];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7544_o = n7543_o;
      13'b0100000000000: n7544_o = n7543_o;
      13'b0010000000000: n7544_o = n7543_o;
      13'b0001000000000: n7544_o = n7543_o;
      13'b0000100000000: n7544_o = n7543_o;
      13'b0000010000000: n7544_o = n7543_o;
      13'b0000001000000: n7544_o = n7543_o;
      13'b0000000100000: n7544_o = n7543_o;
      13'b0000000010000: n7544_o = n7543_o;
      13'b0000000001000: n7544_o = n7543_o;
      13'b0000000000100: n7544_o = n5651_o;
      13'b0000000000010: n7544_o = n7543_o;
      13'b0000000000001: n7544_o = n7543_o;
      default: n7544_o = n7543_o;
    endcase
  assign n7545_o = n1909_o[37];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7546_o = n7545_o;
      13'b0100000000000: n7546_o = n7545_o;
      13'b0010000000000: n7546_o = n7545_o;
      13'b0001000000000: n7546_o = n7545_o;
      13'b0000100000000: n7546_o = n7545_o;
      13'b0000010000000: n7546_o = n7545_o;
      13'b0000001000000: n7546_o = n7545_o;
      13'b0000000100000: n7546_o = n7545_o;
      13'b0000000010000: n7546_o = n7545_o;
      13'b0000000001000: n7546_o = n7545_o;
      13'b0000000000100: n7546_o = n7545_o;
      13'b0000000000010: n7546_o = n7545_o;
      13'b0000000000001: n7546_o = n3106_o;
      default: n7546_o = n7545_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7547_o = n2007_o;
      13'b0100000000000: n7547_o = n2007_o;
      13'b0010000000000: n7547_o = n2007_o;
      13'b0001000000000: n7547_o = n6653_o;
      13'b0000100000000: n7547_o = n2007_o;
      13'b0000010000000: n7547_o = n2007_o;
      13'b0000001000000: n7547_o = n2007_o;
      13'b0000000100000: n7547_o = n2007_o;
      13'b0000000010000: n7547_o = n2007_o;
      13'b0000000001000: n7547_o = n2007_o;
      13'b0000000000100: n7547_o = n2007_o;
      13'b0000000000010: n7547_o = n2007_o;
      13'b0000000000001: n7547_o = n2007_o;
      default: n7547_o = n2007_o;
    endcase
  assign n7548_o = n1909_o[39];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7549_o = n7548_o;
      13'b0100000000000: n7549_o = n7548_o;
      13'b0010000000000: n7549_o = n7548_o;
      13'b0001000000000: n7549_o = n7548_o;
      13'b0000100000000: n7549_o = n7548_o;
      13'b0000010000000: n7549_o = n7548_o;
      13'b0000001000000: n7549_o = n7548_o;
      13'b0000000100000: n7549_o = n7548_o;
      13'b0000000010000: n7549_o = n7548_o;
      13'b0000000001000: n7549_o = n7548_o;
      13'b0000000000100: n7549_o = n7548_o;
      13'b0000000000010: n7549_o = n7548_o;
      13'b0000000000001: n7549_o = n3108_o;
      default: n7549_o = n7548_o;
    endcase
  assign n7550_o = n1909_o[40];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7551_o = n7550_o;
      13'b0100000000000: n7551_o = n7550_o;
      13'b0010000000000: n7551_o = n7550_o;
      13'b0001000000000: n7551_o = n7550_o;
      13'b0000100000000: n7551_o = n7550_o;
      13'b0000010000000: n7551_o = n7550_o;
      13'b0000001000000: n7551_o = n7550_o;
      13'b0000000100000: n7551_o = n7550_o;
      13'b0000000010000: n7551_o = n7550_o;
      13'b0000000001000: n7551_o = n7550_o;
      13'b0000000000100: n7551_o = n5653_o;
      13'b0000000000010: n7551_o = n3308_o;
      13'b0000000000001: n7551_o = n7550_o;
      default: n7551_o = n7550_o;
    endcase
  assign n7552_o = n3110_o[0];
  assign n7553_o = n1909_o[42];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7554_o = n7553_o;
      13'b0100000000000: n7554_o = n7298_o;
      13'b0010000000000: n7554_o = n7553_o;
      13'b0001000000000: n7554_o = n7553_o;
      13'b0000100000000: n7554_o = n7553_o;
      13'b0000010000000: n7554_o = n7553_o;
      13'b0000001000000: n7554_o = n7553_o;
      13'b0000000100000: n7554_o = n7553_o;
      13'b0000000010000: n7554_o = n7553_o;
      13'b0000000001000: n7554_o = n7553_o;
      13'b0000000000100: n7554_o = n5655_o;
      13'b0000000000010: n7554_o = n7553_o;
      13'b0000000000001: n7554_o = n7552_o;
      default: n7554_o = n7553_o;
    endcase
  assign n7555_o = n3110_o[1];
  assign n7556_o = n1909_o[43];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7557_o = n7556_o;
      13'b0100000000000: n7557_o = n7556_o;
      13'b0010000000000: n7557_o = n7556_o;
      13'b0001000000000: n7557_o = n7556_o;
      13'b0000100000000: n7557_o = n7556_o;
      13'b0000010000000: n7557_o = n7556_o;
      13'b0000001000000: n7557_o = n7556_o;
      13'b0000000100000: n7557_o = n7556_o;
      13'b0000000010000: n7557_o = n7556_o;
      13'b0000000001000: n7557_o = n7556_o;
      13'b0000000000100: n7557_o = n5657_o;
      13'b0000000000010: n7557_o = n7556_o;
      13'b0000000000001: n7557_o = n7555_o;
      default: n7557_o = n7556_o;
    endcase
  assign n7558_o = n1909_o[44];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7559_o = n7558_o;
      13'b0100000000000: n7559_o = n7558_o;
      13'b0010000000000: n7559_o = n7558_o;
      13'b0001000000000: n7559_o = n7558_o;
      13'b0000100000000: n7559_o = n7558_o;
      13'b0000010000000: n7559_o = n7558_o;
      13'b0000001000000: n7559_o = n6320_o;
      13'b0000000100000: n7559_o = n7558_o;
      13'b0000000010000: n7559_o = n7558_o;
      13'b0000000001000: n7559_o = n7558_o;
      13'b0000000000100: n7559_o = n5659_o;
      13'b0000000000010: n7559_o = n7558_o;
      13'b0000000000001: n7559_o = n7558_o;
      default: n7559_o = n7558_o;
    endcase
  assign n7560_o = n3309_o[0];
  assign n7561_o = n5663_o[0];
  assign n7562_o = n2162_o[0];
  assign n7563_o = n1909_o[46];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n7564_o = n2037_o ? n7562_o : n7563_o;
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7565_o = n7564_o;
      13'b0100000000000: n7565_o = n7564_o;
      13'b0010000000000: n7565_o = n7564_o;
      13'b0001000000000: n7565_o = n6657_o;
      13'b0000100000000: n7565_o = n7564_o;
      13'b0000010000000: n7565_o = n7564_o;
      13'b0000001000000: n7565_o = n7564_o;
      13'b0000000100000: n7565_o = n7564_o;
      13'b0000000010000: n7565_o = n7564_o;
      13'b0000000001000: n7565_o = n7564_o;
      13'b0000000000100: n7565_o = n7561_o;
      13'b0000000000010: n7565_o = n7560_o;
      13'b0000000000001: n7565_o = n7564_o;
      default: n7565_o = n7564_o;
    endcase
  assign n7566_o = n3309_o[1];
  assign n7567_o = n5663_o[1];
  assign n7568_o = n2162_o[1];
  assign n7569_o = n1909_o[47];
  /* TG68KdotC_Kernel.vhd:1594:17  */
  assign n7570_o = n2037_o ? n7568_o : n7569_o;
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7571_o = n7570_o;
      13'b0100000000000: n7571_o = n7570_o;
      13'b0010000000000: n7571_o = n7570_o;
      13'b0001000000000: n7571_o = n7570_o;
      13'b0000100000000: n7571_o = n7570_o;
      13'b0000010000000: n7571_o = n7570_o;
      13'b0000001000000: n7571_o = n7570_o;
      13'b0000000100000: n7571_o = n7570_o;
      13'b0000000010000: n7571_o = n5990_o;
      13'b0000000001000: n7571_o = n7570_o;
      13'b0000000000100: n7571_o = n7567_o;
      13'b0000000000010: n7571_o = n7566_o;
      13'b0000000000001: n7571_o = n7570_o;
      default: n7571_o = n7570_o;
    endcase
  assign n7572_o = n5663_o[2];
  assign n7573_o = n1909_o[48];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7574_o = n7573_o;
      13'b0100000000000: n7574_o = n7573_o;
      13'b0010000000000: n7574_o = n7573_o;
      13'b0001000000000: n7574_o = n7573_o;
      13'b0000100000000: n7574_o = n7573_o;
      13'b0000010000000: n7574_o = n7573_o;
      13'b0000001000000: n7574_o = n7573_o;
      13'b0000000100000: n7574_o = n7573_o;
      13'b0000000010000: n7574_o = n7573_o;
      13'b0000000001000: n7574_o = n7573_o;
      13'b0000000000100: n7574_o = n7572_o;
      13'b0000000000010: n7574_o = n7573_o;
      13'b0000000000001: n7574_o = n7573_o;
      default: n7574_o = n7573_o;
    endcase
  assign n7575_o = n3341_o[0];
  assign n7576_o = n1909_o[49];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7577_o = n7576_o;
      13'b0100000000000: n7577_o = n7576_o;
      13'b0010000000000: n7577_o = n7576_o;
      13'b0001000000000: n7577_o = n7576_o;
      13'b0000100000000: n7577_o = n7576_o;
      13'b0000010000000: n7577_o = n6420_o;
      13'b0000001000000: n7577_o = n6322_o;
      13'b0000000100000: n7577_o = n7576_o;
      13'b0000000010000: n7577_o = n7576_o;
      13'b0000000001000: n7577_o = n5917_o;
      13'b0000000000100: n7577_o = n5665_o;
      13'b0000000000010: n7577_o = n7575_o;
      13'b0000000000001: n7577_o = n3112_o;
      default: n7577_o = n7576_o;
    endcase
  assign n7578_o = n3341_o[1];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7579_o = n2168_o;
      13'b0100000000000: n7579_o = n2168_o;
      13'b0010000000000: n7579_o = n2168_o;
      13'b0001000000000: n7579_o = n6658_o;
      13'b0000100000000: n7579_o = n2168_o;
      13'b0000010000000: n7579_o = n2168_o;
      13'b0000001000000: n7579_o = n2168_o;
      13'b0000000100000: n7579_o = n2168_o;
      13'b0000000010000: n7579_o = n2168_o;
      13'b0000000001000: n7579_o = n2168_o;
      13'b0000000000100: n7579_o = n2168_o;
      13'b0000000000010: n7579_o = n7578_o;
      13'b0000000000001: n7579_o = n3114_o;
      default: n7579_o = n2168_o;
    endcase
  assign n7580_o = n5668_o[1:0];
  assign n7581_o = n1909_o[52:51];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7582_o = n7581_o;
      13'b0100000000000: n7582_o = n7581_o;
      13'b0010000000000: n7582_o = n7581_o;
      13'b0001000000000: n7582_o = n7581_o;
      13'b0000100000000: n7582_o = n7581_o;
      13'b0000010000000: n7582_o = n7581_o;
      13'b0000001000000: n7582_o = n7581_o;
      13'b0000000100000: n7582_o = n7581_o;
      13'b0000000010000: n7582_o = n7581_o;
      13'b0000000001000: n7582_o = n7581_o;
      13'b0000000000100: n7582_o = n7580_o;
      13'b0000000000010: n7582_o = n7581_o;
      13'b0000000000001: n7582_o = n3116_o;
      default: n7582_o = n7581_o;
    endcase
  assign n7583_o = n5668_o[2];
  assign n7584_o = n1909_o[53];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7585_o = n7584_o;
      13'b0100000000000: n7585_o = n7584_o;
      13'b0010000000000: n7585_o = n7584_o;
      13'b0001000000000: n7585_o = n7584_o;
      13'b0000100000000: n7585_o = n7584_o;
      13'b0000010000000: n7585_o = n7584_o;
      13'b0000001000000: n7585_o = n7584_o;
      13'b0000000100000: n7585_o = n7584_o;
      13'b0000000010000: n7585_o = n7584_o;
      13'b0000000001000: n7585_o = n5724_o;
      13'b0000000000100: n7585_o = n7583_o;
      13'b0000000000010: n7585_o = n7584_o;
      13'b0000000000001: n7585_o = n7584_o;
      default: n7585_o = n7584_o;
    endcase
  assign n7586_o = n5668_o[3];
  assign n7587_o = n1909_o[54];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7588_o = n7587_o;
      13'b0100000000000: n7588_o = n7587_o;
      13'b0010000000000: n7588_o = n7587_o;
      13'b0001000000000: n7588_o = n7587_o;
      13'b0000100000000: n7588_o = n7587_o;
      13'b0000010000000: n7588_o = n7587_o;
      13'b0000001000000: n7588_o = n7587_o;
      13'b0000000100000: n7588_o = n7587_o;
      13'b0000000010000: n7588_o = n7587_o;
      13'b0000000001000: n7588_o = n7587_o;
      13'b0000000000100: n7588_o = n7586_o;
      13'b0000000000010: n7588_o = n7587_o;
      13'b0000000000001: n7588_o = n7587_o;
      default: n7588_o = n7587_o;
    endcase
  assign n7589_o = n3118_o[0];
  assign n7590_o = n5668_o[4];
  assign n7591_o = n1909_o[55];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7592_o = n7591_o;
      13'b0100000000000: n7592_o = n7300_o;
      13'b0010000000000: n7592_o = n7591_o;
      13'b0001000000000: n7592_o = n7591_o;
      13'b0000100000000: n7592_o = n7591_o;
      13'b0000010000000: n7592_o = n7591_o;
      13'b0000001000000: n7592_o = n7591_o;
      13'b0000000100000: n7592_o = n7591_o;
      13'b0000000010000: n7592_o = n7591_o;
      13'b0000000001000: n7592_o = n7591_o;
      13'b0000000000100: n7592_o = n7590_o;
      13'b0000000000010: n7592_o = n7591_o;
      13'b0000000000001: n7592_o = n7589_o;
      default: n7592_o = n7591_o;
    endcase
  assign n7593_o = n3118_o[1];
  assign n7594_o = n1909_o[56];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7595_o = n7594_o;
      13'b0100000000000: n7595_o = n7594_o;
      13'b0010000000000: n7595_o = n7594_o;
      13'b0001000000000: n7595_o = n6659_o;
      13'b0000100000000: n7595_o = n7594_o;
      13'b0000010000000: n7595_o = n6374_o;
      13'b0000001000000: n7595_o = n6324_o;
      13'b0000000100000: n7595_o = n7594_o;
      13'b0000000010000: n7595_o = n7594_o;
      13'b0000000001000: n7595_o = n5921_o;
      13'b0000000000100: n7595_o = n5670_o;
      13'b0000000000010: n7595_o = n7594_o;
      13'b0000000000001: n7595_o = n7593_o;
      default: n7595_o = n7594_o;
    endcase
  assign n7596_o = n1909_o[60:57];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7597_o = n7596_o;
      13'b0100000000000: n7597_o = n7596_o;
      13'b0010000000000: n7597_o = n7596_o;
      13'b0001000000000: n7597_o = n7596_o;
      13'b0000100000000: n7597_o = n7596_o;
      13'b0000010000000: n7597_o = n7596_o;
      13'b0000001000000: n7597_o = n7596_o;
      13'b0000000100000: n7597_o = n7596_o;
      13'b0000000010000: n7597_o = n7596_o;
      13'b0000000001000: n7597_o = n7596_o;
      13'b0000000000100: n7597_o = n5673_o;
      13'b0000000000010: n7597_o = n7596_o;
      13'b0000000000001: n7597_o = n7596_o;
      default: n7597_o = n7596_o;
    endcase
  assign n7598_o = n1909_o[61];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7599_o = n7598_o;
      13'b0100000000000: n7599_o = n7598_o;
      13'b0010000000000: n7599_o = n6920_o;
      13'b0001000000000: n7599_o = n7598_o;
      13'b0000100000000: n7599_o = n7598_o;
      13'b0000010000000: n7599_o = n7598_o;
      13'b0000001000000: n7599_o = n7598_o;
      13'b0000000100000: n7599_o = n7598_o;
      13'b0000000010000: n7599_o = n7598_o;
      13'b0000000001000: n7599_o = n7598_o;
      13'b0000000000100: n7599_o = n7598_o;
      13'b0000000000010: n7599_o = n7598_o;
      13'b0000000000001: n7599_o = n7598_o;
      default: n7599_o = n7598_o;
    endcase
  assign n7600_o = {n2019_o, n2178_o};
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7601_o = n7600_o;
      13'b0100000000000: n7601_o = n7600_o;
      13'b0010000000000: n7601_o = n7600_o;
      13'b0001000000000: n7601_o = n7600_o;
      13'b0000100000000: n7601_o = n7600_o;
      13'b0000010000000: n7601_o = n7600_o;
      13'b0000001000000: n7601_o = n7600_o;
      13'b0000000100000: n7601_o = n7600_o;
      13'b0000000010000: n7601_o = n7600_o;
      13'b0000000001000: n7601_o = n7600_o;
      13'b0000000000100: n7601_o = n5675_o;
      13'b0000000000010: n7601_o = n7600_o;
      13'b0000000000001: n7601_o = n7600_o;
      default: n7601_o = n7600_o;
    endcase
  assign n7602_o = n1909_o[69];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7603_o = n7602_o;
      13'b0100000000000: n7603_o = n7602_o;
      13'b0010000000000: n7603_o = n7602_o;
      13'b0001000000000: n7603_o = n7602_o;
      13'b0000100000000: n7603_o = n7602_o;
      13'b0000010000000: n7603_o = n7602_o;
      13'b0000001000000: n7603_o = n7602_o;
      13'b0000000100000: n7603_o = n7602_o;
      13'b0000000010000: n7603_o = n7602_o;
      13'b0000000001000: n7603_o = n7602_o;
      13'b0000000000100: n7603_o = n5677_o;
      13'b0000000000010: n7603_o = n7602_o;
      13'b0000000000001: n7603_o = n7602_o;
      default: n7603_o = n7602_o;
    endcase
  assign n7604_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7605_o = n7604_o;
      13'b0100000000000: n7605_o = n7302_o;
      13'b0010000000000: n7605_o = n7604_o;
      13'b0001000000000: n7605_o = n7604_o;
      13'b0000100000000: n7605_o = n7604_o;
      13'b0000010000000: n7605_o = n7604_o;
      13'b0000001000000: n7605_o = n7604_o;
      13'b0000000100000: n7605_o = n7604_o;
      13'b0000000010000: n7605_o = n7604_o;
      13'b0000000001000: n7605_o = n7604_o;
      13'b0000000000100: n7605_o = n5679_o;
      13'b0000000000010: n7605_o = n7604_o;
      13'b0000000000001: n7605_o = n3120_o;
      default: n7605_o = n7604_o;
    endcase
  assign n7606_o = n5682_o[0];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7607_o = n2171_o;
      13'b0100000000000: n7607_o = n2171_o;
      13'b0010000000000: n7607_o = n2171_o;
      13'b0001000000000: n7607_o = n2171_o;
      13'b0000100000000: n7607_o = n2171_o;
      13'b0000010000000: n7607_o = n2171_o;
      13'b0000001000000: n7607_o = n2171_o;
      13'b0000000100000: n7607_o = n2171_o;
      13'b0000000010000: n7607_o = n5991_o;
      13'b0000000001000: n7607_o = n5922_o;
      13'b0000000000100: n7607_o = n7606_o;
      13'b0000000000010: n7607_o = n3311_o;
      13'b0000000000001: n7607_o = n3121_o;
      default: n7607_o = n2171_o;
    endcase
  assign n7608_o = n5682_o[1];
  assign n7609_o = n1909_o[74];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7610_o = n7609_o;
      13'b0100000000000: n7610_o = n7609_o;
      13'b0010000000000: n7610_o = n7609_o;
      13'b0001000000000: n7610_o = n7609_o;
      13'b0000100000000: n7610_o = n7609_o;
      13'b0000010000000: n7610_o = n7609_o;
      13'b0000001000000: n7610_o = n7609_o;
      13'b0000000100000: n7610_o = n7609_o;
      13'b0000000010000: n7610_o = n7609_o;
      13'b0000000001000: n7610_o = n7609_o;
      13'b0000000000100: n7610_o = n7608_o;
      13'b0000000000010: n7610_o = n7609_o;
      13'b0000000000001: n7610_o = n7609_o;
      default: n7610_o = n7609_o;
    endcase
  assign n7611_o = n1909_o[80];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7612_o = n7611_o;
      13'b0100000000000: n7612_o = n7611_o;
      13'b0010000000000: n7612_o = n7611_o;
      13'b0001000000000: n7612_o = n7611_o;
      13'b0000100000000: n7612_o = n7611_o;
      13'b0000010000000: n7612_o = n7611_o;
      13'b0000001000000: n7612_o = n6326_o;
      13'b0000000100000: n7612_o = n7611_o;
      13'b0000000010000: n7612_o = n7611_o;
      13'b0000000001000: n7612_o = n7611_o;
      13'b0000000000100: n7612_o = n7611_o;
      13'b0000000000010: n7612_o = n7611_o;
      13'b0000000000001: n7612_o = n7611_o;
      default: n7612_o = n7611_o;
    endcase
  assign n7613_o = n1909_o[82];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7614_o = n7613_o;
      13'b0100000000000: n7614_o = n7613_o;
      13'b0010000000000: n7614_o = n7613_o;
      13'b0001000000000: n7614_o = n7613_o;
      13'b0000100000000: n7614_o = n7613_o;
      13'b0000010000000: n7614_o = n7613_o;
      13'b0000001000000: n7614_o = n7613_o;
      13'b0000000100000: n7614_o = n7613_o;
      13'b0000000010000: n7614_o = n7613_o;
      13'b0000000001000: n7614_o = n7613_o;
      13'b0000000000100: n7614_o = n7613_o;
      13'b0000000000010: n7614_o = n7613_o;
      13'b0000000000001: n7614_o = n3123_o;
      default: n7614_o = n7613_o;
    endcase
  assign n7615_o = n1909_o[84];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7616_o = n7615_o;
      13'b0100000000000: n7616_o = n7615_o;
      13'b0010000000000: n7616_o = n7615_o;
      13'b0001000000000: n7616_o = n7615_o;
      13'b0000100000000: n7616_o = n7615_o;
      13'b0000010000000: n7616_o = n7615_o;
      13'b0000001000000: n7616_o = n7615_o;
      13'b0000000100000: n7616_o = n7615_o;
      13'b0000000010000: n7616_o = n7615_o;
      13'b0000000001000: n7616_o = n7615_o;
      13'b0000000000100: n7616_o = n7615_o;
      13'b0000000000010: n7616_o = n7615_o;
      13'b0000000000001: n7616_o = n3125_o;
      default: n7616_o = n7615_o;
    endcase
  assign n7617_o = n1909_o[85];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7618_o = n7617_o;
      13'b0100000000000: n7618_o = n7617_o;
      13'b0010000000000: n7618_o = n6922_o;
      13'b0001000000000: n7618_o = n7617_o;
      13'b0000100000000: n7618_o = n7617_o;
      13'b0000010000000: n7618_o = n7617_o;
      13'b0000001000000: n7618_o = n7617_o;
      13'b0000000100000: n7618_o = n7617_o;
      13'b0000000010000: n7618_o = n7617_o;
      13'b0000000001000: n7618_o = n7617_o;
      13'b0000000000100: n7618_o = n7617_o;
      13'b0000000000010: n7618_o = n7617_o;
      13'b0000000000001: n7618_o = n7617_o;
      default: n7618_o = n7617_o;
    endcase
  assign n7619_o = n1909_o[86];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7620_o = n7619_o;
      13'b0100000000000: n7620_o = n7619_o;
      13'b0010000000000: n7620_o = n7619_o;
      13'b0001000000000: n7620_o = n7619_o;
      13'b0000100000000: n7620_o = n7619_o;
      13'b0000010000000: n7620_o = n7619_o;
      13'b0000001000000: n7620_o = n7619_o;
      13'b0000000100000: n7620_o = n7619_o;
      13'b0000000010000: n7620_o = n7619_o;
      13'b0000000001000: n7620_o = n7619_o;
      13'b0000000000100: n7620_o = n7619_o;
      13'b0000000000010: n7620_o = n7619_o;
      13'b0000000000001: n7620_o = n3127_o;
      default: n7620_o = n7619_o;
    endcase
  assign n7621_o = n6013_o[0];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7623_o = 1'b0;
      13'b0100000000000: n7623_o = 1'b0;
      13'b0010000000000: n7623_o = 1'b0;
      13'b0001000000000: n7623_o = 1'b0;
      13'b0000100000000: n7623_o = 1'b0;
      13'b0000010000000: n7623_o = 1'b0;
      13'b0000001000000: n7623_o = 1'b0;
      13'b0000000100000: n7623_o = n7621_o;
      13'b0000000010000: n7623_o = 1'b0;
      13'b0000000001000: n7623_o = 1'b0;
      13'b0000000000100: n7623_o = n5686_o;
      13'b0000000000010: n7623_o = n3344_o;
      13'b0000000000001: n7623_o = n3129_o;
      default: n7623_o = 1'b0;
    endcase
  assign n7624_o = n6013_o[1];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7626_o = 1'b0;
      13'b0100000000000: n7626_o = 1'b0;
      13'b0010000000000: n7626_o = 1'b0;
      13'b0001000000000: n7626_o = 1'b0;
      13'b0000100000000: n7626_o = 1'b0;
      13'b0000010000000: n7626_o = 1'b0;
      13'b0000001000000: n7626_o = 1'b0;
      13'b0000000100000: n7626_o = n7624_o;
      13'b0000000010000: n7626_o = 1'b0;
      13'b0000000001000: n7626_o = 1'b0;
      13'b0000000000100: n7626_o = 1'b0;
      13'b0000000000010: n7626_o = 1'b0;
      13'b0000000000001: n7626_o = 1'b0;
      default: n7626_o = 1'b0;
    endcase
  assign n7627_o = n5688_o[0];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7629_o = 1'b0;
      13'b0100000000000: n7629_o = 1'b0;
      13'b0010000000000: n7629_o = 1'b0;
      13'b0001000000000: n7629_o = 1'b0;
      13'b0000100000000: n7629_o = 1'b0;
      13'b0000010000000: n7629_o = 1'b0;
      13'b0000001000000: n7629_o = 1'b0;
      13'b0000000100000: n7629_o = 1'b0;
      13'b0000000010000: n7629_o = 1'b0;
      13'b0000000001000: n7629_o = 1'b0;
      13'b0000000000100: n7629_o = n7627_o;
      13'b0000000000010: n7629_o = 1'b0;
      13'b0000000000001: n7629_o = 1'b0;
      default: n7629_o = 1'b0;
    endcase
  assign n7630_o = n5688_o[1];
  assign n7631_o = n5924_o[0];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7633_o = 1'b0;
      13'b0100000000000: n7633_o = 1'b0;
      13'b0010000000000: n7633_o = n6924_o;
      13'b0001000000000: n7633_o = 1'b0;
      13'b0000100000000: n7633_o = 1'b0;
      13'b0000010000000: n7633_o = n6450_o;
      13'b0000001000000: n7633_o = n6328_o;
      13'b0000000100000: n7633_o = 1'b0;
      13'b0000000010000: n7633_o = 1'b0;
      13'b0000000001000: n7633_o = n7631_o;
      13'b0000000000100: n7633_o = n7630_o;
      13'b0000000000010: n7633_o = 1'b0;
      13'b0000000000001: n7633_o = n3131_o;
      default: n7633_o = 1'b0;
    endcase
  assign n7634_o = n5924_o[1];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7636_o = 1'b0;
      13'b0100000000000: n7636_o = 1'b0;
      13'b0010000000000: n7636_o = 1'b0;
      13'b0001000000000: n7636_o = 1'b0;
      13'b0000100000000: n7636_o = 1'b0;
      13'b0000010000000: n7636_o = 1'b0;
      13'b0000001000000: n7636_o = 1'b0;
      13'b0000000100000: n7636_o = 1'b0;
      13'b0000000010000: n7636_o = 1'b0;
      13'b0000000001000: n7636_o = n7634_o;
      13'b0000000000100: n7636_o = 1'b0;
      13'b0000000000010: n7636_o = 1'b0;
      13'b0000000000001: n7636_o = 1'b0;
      default: n7636_o = 1'b0;
    endcase
  assign n7637_o = n3133_o[0];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7639_o = 1'b0;
      13'b0100000000000: n7639_o = 1'b0;
      13'b0010000000000: n7639_o = 1'b0;
      13'b0001000000000: n7639_o = 1'b0;
      13'b0000100000000: n7639_o = 1'b0;
      13'b0000010000000: n7639_o = 1'b0;
      13'b0000001000000: n7639_o = n6330_o;
      13'b0000000100000: n7639_o = 1'b0;
      13'b0000000010000: n7639_o = 1'b0;
      13'b0000000001000: n7639_o = 1'b0;
      13'b0000000000100: n7639_o = 1'b0;
      13'b0000000000010: n7639_o = 1'b0;
      13'b0000000000001: n7639_o = n7637_o;
      default: n7639_o = 1'b0;
    endcase
  assign n7640_o = n3133_o[1];
  assign n7641_o = n5690_o[0];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7643_o = 1'b0;
      13'b0100000000000: n7643_o = 1'b0;
      13'b0010000000000: n7643_o = n6926_o;
      13'b0001000000000: n7643_o = 1'b0;
      13'b0000100000000: n7643_o = 1'b0;
      13'b0000010000000: n7643_o = 1'b0;
      13'b0000001000000: n7643_o = 1'b0;
      13'b0000000100000: n7643_o = 1'b0;
      13'b0000000010000: n7643_o = 1'b0;
      13'b0000000001000: n7643_o = 1'b0;
      13'b0000000000100: n7643_o = n7641_o;
      13'b0000000000010: n7643_o = 1'b0;
      13'b0000000000001: n7643_o = n7640_o;
      default: n7643_o = 1'b0;
    endcase
  assign n7644_o = n3133_o[2];
  assign n7645_o = n5690_o[1];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7647_o = 1'b0;
      13'b0100000000000: n7647_o = 1'b0;
      13'b0010000000000: n7647_o = 1'b0;
      13'b0001000000000: n7647_o = n6663_o;
      13'b0000100000000: n7647_o = 1'b0;
      13'b0000010000000: n7647_o = 1'b0;
      13'b0000001000000: n7647_o = 1'b0;
      13'b0000000100000: n7647_o = 1'b0;
      13'b0000000010000: n7647_o = 1'b0;
      13'b0000000001000: n7647_o = 1'b0;
      13'b0000000000100: n7647_o = n7645_o;
      13'b0000000000010: n7647_o = 1'b0;
      13'b0000000000001: n7647_o = n7644_o;
      default: n7647_o = 1'b0;
    endcase
  assign n7648_o = n3133_o[3];
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7650_o = 1'b0;
      13'b0100000000000: n7650_o = 1'b0;
      13'b0010000000000: n7650_o = 1'b0;
      13'b0001000000000: n7650_o = n6665_o;
      13'b0000100000000: n7650_o = 1'b0;
      13'b0000010000000: n7650_o = 1'b0;
      13'b0000001000000: n7650_o = 1'b0;
      13'b0000000100000: n7650_o = 1'b0;
      13'b0000000010000: n7650_o = 1'b0;
      13'b0000000001000: n7650_o = 1'b0;
      13'b0000000000100: n7650_o = 1'b0;
      13'b0000000000010: n7650_o = 1'b0;
      13'b0000000000001: n7650_o = n7648_o;
      default: n7650_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7652_o = 1'b0;
      13'b0100000000000: n7652_o = n7303_o;
      13'b0010000000000: n7652_o = 1'b0;
      13'b0001000000000: n7652_o = 1'b0;
      13'b0000100000000: n7652_o = 1'b0;
      13'b0000010000000: n7652_o = 1'b0;
      13'b0000001000000: n7652_o = 1'b0;
      13'b0000000100000: n7652_o = 1'b0;
      13'b0000000010000: n7652_o = 1'b0;
      13'b0000000001000: n7652_o = 1'b0;
      13'b0000000000100: n7652_o = 1'b0;
      13'b0000000000010: n7652_o = 1'b0;
      13'b0000000000001: n7652_o = 1'b0;
      default: n7652_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7654_o = 1'b0;
      13'b0100000000000: n7654_o = 1'b0;
      13'b0010000000000: n7654_o = 1'b0;
      13'b0001000000000: n7654_o = n6667_o;
      13'b0000100000000: n7654_o = 1'b0;
      13'b0000010000000: n7654_o = 1'b0;
      13'b0000001000000: n7654_o = 1'b0;
      13'b0000000100000: n7654_o = 1'b0;
      13'b0000000010000: n7654_o = 1'b0;
      13'b0000000001000: n7654_o = 1'b0;
      13'b0000000000100: n7654_o = 1'b0;
      13'b0000000000010: n7654_o = 1'b0;
      13'b0000000000001: n7654_o = 1'b0;
      default: n7654_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7656_o = 1'b0;
      13'b0100000000000: n7656_o = 1'b0;
      13'b0010000000000: n7656_o = 1'b0;
      13'b0001000000000: n7656_o = 1'b0;
      13'b0000100000000: n7656_o = 1'b0;
      13'b0000010000000: n7656_o = 1'b0;
      13'b0000001000000: n7656_o = 1'b0;
      13'b0000000100000: n7656_o = 1'b0;
      13'b0000000010000: n7656_o = 1'b0;
      13'b0000000001000: n7656_o = 1'b0;
      13'b0000000000100: n7656_o = n5691_o;
      13'b0000000000010: n7656_o = 1'b0;
      13'b0000000000001: n7656_o = 1'b0;
      default: n7656_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7658_o = 1'b0;
      13'b0100000000000: n7658_o = 1'b0;
      13'b0010000000000: n7658_o = n6928_o;
      13'b0001000000000: n7658_o = 1'b0;
      13'b0000100000000: n7658_o = 1'b0;
      13'b0000010000000: n7658_o = 1'b0;
      13'b0000001000000: n7658_o = 1'b0;
      13'b0000000100000: n7658_o = 1'b0;
      13'b0000000010000: n7658_o = 1'b0;
      13'b0000000001000: n7658_o = 1'b0;
      13'b0000000000100: n7658_o = 1'b0;
      13'b0000000000010: n7658_o = 1'b0;
      13'b0000000000001: n7658_o = 1'b0;
      default: n7658_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7660_o = 1'b0;
      13'b0100000000000: n7660_o = 1'b0;
      13'b0010000000000: n7660_o = 1'b0;
      13'b0001000000000: n7660_o = 1'b0;
      13'b0000100000000: n7660_o = 1'b0;
      13'b0000010000000: n7660_o = 1'b0;
      13'b0000001000000: n7660_o = n6332_o;
      13'b0000000100000: n7660_o = 1'b0;
      13'b0000000010000: n7660_o = 1'b0;
      13'b0000000001000: n7660_o = 1'b0;
      13'b0000000000100: n7660_o = n5693_o;
      13'b0000000000010: n7660_o = 1'b0;
      13'b0000000000001: n7660_o = 1'b0;
      default: n7660_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7662_o = 1'b0;
      13'b0100000000000: n7662_o = 1'b0;
      13'b0010000000000: n7662_o = 1'b0;
      13'b0001000000000: n7662_o = 1'b0;
      13'b0000100000000: n7662_o = 1'b0;
      13'b0000010000000: n7662_o = 1'b0;
      13'b0000001000000: n7662_o = 1'b0;
      13'b0000000100000: n7662_o = 1'b0;
      13'b0000000010000: n7662_o = 1'b0;
      13'b0000000001000: n7662_o = 1'b0;
      13'b0000000000100: n7662_o = 1'b0;
      13'b0000000000010: n7662_o = 1'b0;
      13'b0000000000001: n7662_o = n3135_o;
      default: n7662_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7664_o = 1'b0;
      13'b0100000000000: n7664_o = 1'b0;
      13'b0010000000000: n7664_o = 1'b0;
      13'b0001000000000: n7664_o = 1'b0;
      13'b0000100000000: n7664_o = 1'b0;
      13'b0000010000000: n7664_o = 1'b0;
      13'b0000001000000: n7664_o = 1'b0;
      13'b0000000100000: n7664_o = 1'b0;
      13'b0000000010000: n7664_o = 1'b0;
      13'b0000000001000: n7664_o = 1'b0;
      13'b0000000000100: n7664_o = n5695_o;
      13'b0000000000010: n7664_o = 1'b0;
      13'b0000000000001: n7664_o = 1'b0;
      default: n7664_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7666_o = 1'b0;
      13'b0100000000000: n7666_o = 1'b0;
      13'b0010000000000: n7666_o = 1'b0;
      13'b0001000000000: n7666_o = 1'b0;
      13'b0000100000000: n7666_o = 1'b0;
      13'b0000010000000: n7666_o = 1'b0;
      13'b0000001000000: n7666_o = 1'b0;
      13'b0000000100000: n7666_o = 1'b0;
      13'b0000000010000: n7666_o = 1'b0;
      13'b0000000001000: n7666_o = n5926_o;
      13'b0000000000100: n7666_o = 1'b0;
      13'b0000000000010: n7666_o = 1'b0;
      13'b0000000000001: n7666_o = 1'b0;
      default: n7666_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7668_o = 1'b0;
      13'b0100000000000: n7668_o = n7305_o;
      13'b0010000000000: n7668_o = 1'b0;
      13'b0001000000000: n7668_o = n6669_o;
      13'b0000100000000: n7668_o = 1'b0;
      13'b0000010000000: n7668_o = 1'b0;
      13'b0000001000000: n7668_o = n6334_o;
      13'b0000000100000: n7668_o = 1'b0;
      13'b0000000010000: n7668_o = 1'b0;
      13'b0000000001000: n7668_o = n5928_o;
      13'b0000000000100: n7668_o = n5697_o;
      13'b0000000000010: n7668_o = 1'b0;
      13'b0000000000001: n7668_o = n3137_o;
      default: n7668_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7670_o = 1'b0;
      13'b0100000000000: n7670_o = 1'b0;
      13'b0010000000000: n7670_o = 1'b0;
      13'b0001000000000: n7670_o = 1'b0;
      13'b0000100000000: n7670_o = 1'b0;
      13'b0000010000000: n7670_o = 1'b0;
      13'b0000001000000: n7670_o = 1'b0;
      13'b0000000100000: n7670_o = 1'b0;
      13'b0000000010000: n7670_o = 1'b0;
      13'b0000000001000: n7670_o = 1'b0;
      13'b0000000000100: n7670_o = n5699_o;
      13'b0000000000010: n7670_o = 1'b0;
      13'b0000000000001: n7670_o = 1'b0;
      default: n7670_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7672_o = 1'b0;
      13'b0100000000000: n7672_o = 1'b0;
      13'b0010000000000: n7672_o = 1'b0;
      13'b0001000000000: n7672_o = 1'b0;
      13'b0000100000000: n7672_o = 1'b0;
      13'b0000010000000: n7672_o = 1'b0;
      13'b0000001000000: n7672_o = 1'b0;
      13'b0000000100000: n7672_o = 1'b0;
      13'b0000000010000: n7672_o = 1'b0;
      13'b0000000001000: n7672_o = 1'b0;
      13'b0000000000100: n7672_o = n5701_o;
      13'b0000000000010: n7672_o = 1'b0;
      13'b0000000000001: n7672_o = 1'b0;
      default: n7672_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7674_o = 1'b0;
      13'b0100000000000: n7674_o = 1'b0;
      13'b0010000000000: n7674_o = 1'b0;
      13'b0001000000000: n7674_o = 1'b0;
      13'b0000100000000: n7674_o = 1'b0;
      13'b0000010000000: n7674_o = 1'b0;
      13'b0000001000000: n7674_o = 1'b0;
      13'b0000000100000: n7674_o = 1'b0;
      13'b0000000010000: n7674_o = 1'b0;
      13'b0000000001000: n7674_o = 1'b0;
      13'b0000000000100: n7674_o = n5703_o;
      13'b0000000000010: n7674_o = 1'b0;
      13'b0000000000001: n7674_o = 1'b0;
      default: n7674_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7676_o = 2'b00;
      13'b0100000000000: n7676_o = 2'b00;
      13'b0010000000000: n7676_o = 2'b00;
      13'b0001000000000: n7676_o = 2'b00;
      13'b0000100000000: n7676_o = 2'b00;
      13'b0000010000000: n7676_o = 2'b00;
      13'b0000001000000: n7676_o = 2'b00;
      13'b0000000100000: n7676_o = 2'b00;
      13'b0000000010000: n7676_o = 2'b00;
      13'b0000000001000: n7676_o = 2'b00;
      13'b0000000000100: n7676_o = n5706_o;
      13'b0000000000010: n7676_o = 2'b00;
      13'b0000000000001: n7676_o = 2'b00;
      default: n7676_o = 2'b00;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7678_o = 1'b0;
      13'b0100000000000: n7678_o = n7306_o;
      13'b0010000000000: n7678_o = n6930_o;
      13'b0001000000000: n7678_o = 1'b0;
      13'b0000100000000: n7678_o = 1'b0;
      13'b0000010000000: n7678_o = n6452_o;
      13'b0000001000000: n7678_o = n6335_o;
      13'b0000000100000: n7678_o = n6015_o;
      13'b0000000010000: n7678_o = 1'b0;
      13'b0000000001000: n7678_o = n5929_o;
      13'b0000000000100: n7678_o = n5708_o;
      13'b0000000000010: n7678_o = n3346_o;
      13'b0000000000001: n7678_o = n3138_o;
      default: n7678_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7680_o = 2'b00;
      13'b0100000000000: n7680_o = n7308_o;
      13'b0010000000000: n7680_o = 2'b00;
      13'b0001000000000: n7680_o = 2'b00;
      13'b0000100000000: n7680_o = 2'b00;
      13'b0000010000000: n7680_o = 2'b00;
      13'b0000001000000: n7680_o = 2'b00;
      13'b0000000100000: n7680_o = 2'b00;
      13'b0000000010000: n7680_o = 2'b00;
      13'b0000000001000: n7680_o = 2'b00;
      13'b0000000000100: n7680_o = 2'b00;
      13'b0000000000010: n7680_o = 2'b00;
      13'b0000000000001: n7680_o = 2'b00;
      default: n7680_o = 2'b00;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7682_o = 2'b00;
      13'b0100000000000: n7682_o = 2'b00;
      13'b0010000000000: n7682_o = 2'b00;
      13'b0001000000000: n7682_o = 2'b00;
      13'b0000100000000: n7682_o = 2'b00;
      13'b0000010000000: n7682_o = 2'b00;
      13'b0000001000000: n7682_o = n6337_o;
      13'b0000000100000: n7682_o = 2'b00;
      13'b0000000010000: n7682_o = 2'b00;
      13'b0000000001000: n7682_o = 2'b00;
      13'b0000000000100: n7682_o = 2'b00;
      13'b0000000000010: n7682_o = 2'b00;
      13'b0000000000001: n7682_o = 2'b00;
      default: n7682_o = 2'b00;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7684_o = 1'b0;
      13'b0100000000000: n7684_o = 1'b0;
      13'b0010000000000: n7684_o = 1'b0;
      13'b0001000000000: n7684_o = 1'b0;
      13'b0000100000000: n7684_o = 1'b0;
      13'b0000010000000: n7684_o = 1'b0;
      13'b0000001000000: n7684_o = 1'b0;
      13'b0000000100000: n7684_o = 1'b0;
      13'b0000000010000: n7684_o = 1'b0;
      13'b0000000001000: n7684_o = 1'b0;
      13'b0000000000100: n7684_o = n5709_o;
      13'b0000000000010: n7684_o = 1'b0;
      13'b0000000000001: n7684_o = 1'b0;
      default: n7684_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:1653:17  */
  always @*
    case (n7453_o)
      13'b1000000000000: n7685_o = n2180_o;
      13'b0100000000000: n7685_o = n7309_o;
      13'b0010000000000: n7685_o = n6709_o;
      13'b0001000000000: n7685_o = n6670_o;
      13'b0000100000000: n7685_o = n2180_o;
      13'b0000010000000: n7685_o = n2180_o;
      13'b0000001000000: n7685_o = n6338_o;
      13'b0000000100000: n7685_o = n2180_o;
      13'b0000000010000: n7685_o = n5992_o;
      13'b0000000001000: n7685_o = n5930_o;
      13'b0000000000100: n7685_o = n5710_o;
      13'b0000000000010: n7685_o = n3313_o;
      13'b0000000000001: n7685_o = n3139_o;
      default: n7685_o = n2180_o;
    endcase
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7686_o = n2184_o ? make_berr : n7454_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7687_o = n2184_o ? n1921_o : n7456_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7688_o = n2184_o ? datatype : n7457_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7689_o = n2184_o ? n2026_o : n7458_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7690_o = n2184_o ? n2148_o : n7459_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7692_o = n2184_o ? 1'b0 : n7461_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7694_o = n2184_o ? n2151_o : n7462_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7696_o = n2184_o ? 1'b0 : n7464_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7699_o = n2184_o ? 1'b0 : n7466_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7701_o = n2184_o ? n2015_o : n7467_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7703_o = n2184_o ? 1'b0 : n7469_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7706_o = n2184_o ? 1'b0 : n7471_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7709_o = n2184_o ? 1'b0 : n7473_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7712_o = n2184_o ? 1'b0 : n7475_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7715_o = n2184_o ? 1'b0 : n7477_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7718_o = n2184_o ? 1'b0 : n7479_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7721_o = n2184_o ? 1'b0 : n7481_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7724_o = n2184_o ? 1'b0 : n7483_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7727_o = n2184_o ? 1'b0 : n7485_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7730_o = n2184_o ? 1'b0 : n7487_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7732_o = n2184_o ? n1900_o : n7488_o;
  assign n7733_o = {n7498_o, n7493_o};
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7734_o = n2184_o ? n1906_o : n7733_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7736_o = n2184_o ? 1'b0 : n7500_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7738_o = n2184_o ? n2154_o : n7501_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7740_o = n2184_o ? 1'b0 : n7504_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7744_o = n2184_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7747_o = n2184_o ? 1'b0 : n7506_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7750_o = n2184_o ? 1'b0 : n7509_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7753_o = n2184_o ? 1'b0 : n7511_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7756_o = n2184_o ? 1'b0 : n7513_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7759_o = n2184_o ? 1'b0 : n7515_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7762_o = n2184_o ? 1'b1 : n7520_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7765_o = n2184_o ? 1'b0 : n7522_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7768_o = n2184_o ? 1'b0 : n7524_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7771_o = n2184_o ? 1'b0 : n7526_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7774_o = n2184_o ? 1'b0 : n7528_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7777_o = n2184_o ? 1'b0 : n7530_o;
  assign n7779_o = {n7551_o, n7549_o, n7547_o, n7546_o, n7544_o};
  assign n7780_o = {n7559_o, n7557_o, n7554_o};
  assign n7781_o = {n7599_o, n7597_o, n7595_o, n7592_o, n7588_o, n7585_o, n7582_o, n7579_o, n7577_o, n7574_o, n7571_o, n7565_o};
  assign n7782_o = {n7610_o, n7607_o};
  assign n7783_o = {n7620_o, n7618_o, n7616_o};
  assign n7784_o = n1909_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7785_o = n2184_o ? n7784_o : n7532_o;
  assign n7786_o = n1909_o[19:17];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7787_o = n2184_o ? n7786_o : n7534_o;
  assign n7788_o = n1909_o[24];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7789_o = n2184_o ? n7788_o : n7536_o;
  assign n7790_o = n1909_o[26];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7791_o = n2184_o ? n7790_o : n7538_o;
  assign n7792_o = n1909_o[29];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7793_o = n2184_o ? n7792_o : n7540_o;
  assign n7794_o = n1909_o[34];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7795_o = n2184_o ? n7794_o : n7542_o;
  assign n7796_o = n1909_o[37:36];
  assign n7797_o = {n1940_o, n2007_o, n7796_o};
  assign n7799_o = n1909_o[44:42];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7800_o = n2184_o ? n7799_o : n7780_o;
  assign n7801_o = {n2179_o, n2168_o, n2177_o, n2166_o};
  assign n7803_o = {n2019_o, n2178_o};
  assign n7805_o = n1909_o[69];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7806_o = n2184_o ? n7805_o : n7603_o;
  assign n7807_o = n1909_o[71];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7808_o = n2184_o ? n7807_o : n7605_o;
  assign n7809_o = n1909_o[74];
  assign n7810_o = {n7809_o, n2171_o};
  assign n7812_o = n1909_o[80];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7813_o = n2184_o ? n7812_o : n7612_o;
  assign n7814_o = n1909_o[82];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7815_o = n2184_o ? n7814_o : n7614_o;
  assign n7820_o = n1909_o[16:1];
  assign n7821_o = n1909_o[23];
  assign n7826_o = n1909_o[33:30];
  assign n7827_o = n1909_o[35];
  assign n7828_o = n1909_o[45];
  assign n7831_o = n1909_o[72];
  assign n7832_o = n1909_o[70];
  assign n7836_o = n1909_o[81];
  assign n7838_o = {n7666_o, n7664_o, n7662_o, n7660_o, n7658_o, n7656_o, n7654_o, n7652_o, n7650_o, n7647_o, n7643_o, n7639_o, n7636_o, n7633_o, n7629_o, n7626_o, n7623_o};
  assign n7839_o = {n7678_o, n7676_o, n7674_o, n7672_o};
  assign n7840_o = {n7682_o, n7680_o};
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7842_o = n2184_o ? 17'b00000000000000000 : n7838_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7844_o = n2184_o ? 1'b0 : n7668_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7846_o = n2184_o ? 1'b0 : n7670_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7850_o = n2184_o ? 4'b0000 : n7840_o;
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7852_o = n2184_o ? 1'b0 : n7684_o;
  assign n7858_o = n7853_o[27];
  assign n7860_o = n7853_o[29];
  assign n7862_o = n7853_o[74:35];
  assign n7863_o = n7853_o[87:79];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7864_o = n2184_o ? n2180_o : n7685_o;
  /* TG68KdotC_Kernel.vhd:3201:36  */
  assign n7865_o = set_exec[8];
  /* TG68KdotC_Kernel.vhd:3201:44  */
  assign n7866_o = ~n7865_o;
  /* TG68KdotC_Kernel.vhd:3201:60  */
  assign n7867_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:3201:63  */
  assign n7868_o = ~n7867_o;
  /* TG68KdotC_Kernel.vhd:3201:77  */
  assign n7869_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:3201:89  */
  assign n7871_o = n7869_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:3201:68  */
  assign n7872_o = n7868_o | n7871_o;
  /* TG68KdotC_Kernel.vhd:3201:49  */
  assign n7873_o = n7872_o & n7866_o;
  assign n7875_o = n7847_o[4];
  assign n7876_o = n7839_o[4];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7877_o = n2184_o ? n7875_o : n7876_o;
  /* TG68KdotC_Kernel.vhd:3201:25  */
  assign n7878_o = n7873_o ? 1'b1 : n7877_o;
  /* TG68KdotC_Kernel.vhd:3204:34  */
  assign n7879_o = opcode[8];
  /* TG68KdotC_Kernel.vhd:3209:42  */
  assign n7881_o = opcode[3];
  /* TG68KdotC_Kernel.vhd:3209:33  */
  assign n7883_o = n7881_o ? 1'b1 : n7712_o;
  /* TG68KdotC_Kernel.vhd:3212:33  */
  assign n7885_o = setexecopc ? 1'b1 : n7730_o;
  /* TG68KdotC_Kernel.vhd:3199:17  */
  assign n7887_o = n7893_o ? 1'b1 : n7699_o;
  /* TG68KdotC_Kernel.vhd:3204:25  */
  assign n7888_o = n7879_o ? n7712_o : n7883_o;
  /* TG68KdotC_Kernel.vhd:3204:25  */
  assign n7890_o = n7879_o ? n7715_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3204:25  */
  assign n7891_o = n7879_o ? n7730_o : n7885_o;
  /* TG68KdotC_Kernel.vhd:3199:17  */
  assign n7892_o = n7899_o ? 1'b1 : n7844_o;
  /* TG68KdotC_Kernel.vhd:3199:17  */
  assign n7893_o = n7879_o & build_logical;
  /* TG68KdotC_Kernel.vhd:3199:17  */
  assign n7894_o = build_logical ? n7888_o : n7712_o;
  /* TG68KdotC_Kernel.vhd:3199:17  */
  assign n7895_o = build_logical ? n7890_o : n7715_o;
  /* TG68KdotC_Kernel.vhd:3199:17  */
  assign n7896_o = build_logical ? n7891_o : n7730_o;
  /* TG68KdotC_Kernel.vhd:3199:17  */
  assign n7898_o = build_logical ? 1'b1 : n7768_o;
  /* TG68KdotC_Kernel.vhd:3199:17  */
  assign n7899_o = n7879_o & build_logical;
  assign n7900_o = n7847_o[4];
  assign n7901_o = n7839_o[4];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7902_o = n2184_o ? n7900_o : n7901_o;
  /* TG68KdotC_Kernel.vhd:3199:17  */
  assign n7903_o = build_logical ? n7878_o : n7902_o;
  assign n7904_o = n7847_o[3:0];
  assign n7905_o = n7839_o[3:0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7906_o = n2184_o ? n7904_o : n7905_o;
  /* TG68KdotC_Kernel.vhd:3224:34  */
  assign n7909_o = opcode[3];
  /* TG68KdotC_Kernel.vhd:3226:50  */
  assign n7910_o = opcode[2:0];
  /* TG68KdotC_Kernel.vhd:3226:62  */
  assign n7912_o = n7910_o == 3'b111;
  assign n7914_o = n7801_o[4];
  assign n7915_o = n7781_o[4];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7916_o = n2184_o ? n7914_o : n7915_o;
  /* TG68KdotC_Kernel.vhd:3226:41  */
  assign n7917_o = n7912_o ? 1'b1 : n7916_o;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n7921_o = n7957_o ? 2'b10 : n7689_o;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n7923_o = n7962_o ? 1'b1 : n7724_o;
  assign n7924_o = n7797_o[2];
  assign n7925_o = n7779_o[2];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7926_o = n2184_o ? n7924_o : n7925_o;
  /* TG68KdotC_Kernel.vhd:3225:33  */
  assign n7927_o = decodeopc ? 1'b1 : n7926_o;
  assign n7928_o = n7801_o[1];
  assign n7929_o = n7781_o[1];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7930_o = n2184_o ? n7928_o : n7929_o;
  /* TG68KdotC_Kernel.vhd:3225:33  */
  assign n7931_o = decodeopc ? 1'b1 : n7930_o;
  assign n7932_o = n7801_o[4];
  assign n7933_o = n7781_o[4];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7934_o = n2184_o ? n7932_o : n7933_o;
  /* TG68KdotC_Kernel.vhd:3225:33  */
  assign n7935_o = decodeopc ? n7917_o : n7934_o;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n7937_o = n7997_o ? 7'b0100001 : n7864_o;
  /* TG68KdotC_Kernel.vhd:3224:25  */
  assign n7939_o = decodeopc & n7909_o;
  /* TG68KdotC_Kernel.vhd:3224:25  */
  assign n7940_o = decodeopc & n7909_o;
  /* TG68KdotC_Kernel.vhd:3224:25  */
  assign n7942_o = n7909_o ? n7896_o : 1'b1;
  assign n7943_o = n7797_o[2];
  assign n7944_o = n7779_o[2];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7945_o = n2184_o ? n7943_o : n7944_o;
  /* TG68KdotC_Kernel.vhd:3224:25  */
  assign n7946_o = n7909_o ? n7927_o : n7945_o;
  assign n7947_o = n7801_o[1];
  assign n7948_o = n7781_o[1];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7949_o = n2184_o ? n7947_o : n7948_o;
  /* TG68KdotC_Kernel.vhd:3224:25  */
  assign n7950_o = n7909_o ? n7931_o : n7949_o;
  assign n7951_o = n7801_o[4];
  assign n7952_o = n7781_o[4];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7953_o = n2184_o ? n7951_o : n7952_o;
  /* TG68KdotC_Kernel.vhd:3224:25  */
  assign n7954_o = n7909_o ? n7935_o : n7953_o;
  /* TG68KdotC_Kernel.vhd:3224:25  */
  assign n7955_o = n7909_o ? n7903_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3224:25  */
  assign n7956_o = decodeopc & n7909_o;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n7957_o = n7939_o & build_bcd;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n7959_o = build_bcd ? 1'b1 : n7887_o;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n7961_o = build_bcd ? 1'b1 : n7895_o;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n7962_o = n7940_o & build_bcd;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n7963_o = build_bcd ? n7942_o : n7896_o;
  assign n7964_o = n7797_o[2];
  assign n7965_o = n7779_o[2];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7966_o = n2184_o ? n7964_o : n7965_o;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n7967_o = build_bcd ? n7946_o : n7966_o;
  assign n7968_o = n7801_o[1];
  assign n7969_o = n7781_o[1];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7970_o = n2184_o ? n7968_o : n7969_o;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n7971_o = build_bcd ? n7950_o : n7970_o;
  assign n7972_o = n7801_o[4];
  assign n7973_o = n7781_o[4];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7974_o = n2184_o ? n7972_o : n7973_o;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n7975_o = build_bcd ? n7954_o : n7974_o;
  assign n7985_o = n7801_o[0];
  assign n7986_o = n7781_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n7987_o = n2184_o ? n7985_o : n7986_o;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n7994_o = build_bcd ? 1'b1 : n7892_o;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n7995_o = build_bcd ? 1'b1 : n7846_o;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n7996_o = build_bcd ? n7955_o : n7903_o;
  /* TG68KdotC_Kernel.vhd:3219:17  */
  assign n7997_o = n7956_o & build_bcd;
  /* TG68KdotC_Kernel.vhd:3246:33  */
  assign n7998_o = ~trapd;
  /* TG68KdotC_Kernel.vhd:3244:17  */
  assign n8000_o = n8001_o ? 1'b1 : n7703_o;
  /* TG68KdotC_Kernel.vhd:3244:17  */
  assign n8001_o = n7998_o & set_z_error;
  /* TG68KdotC_Kernel.vhd:3244:17  */
  assign n8003_o = set_z_error ? 1'b1 : n7762_o;
  /* TG68KdotC_Kernel.vhd:3257:25  */
  assign n8005_o = clkena_lw ? trapmake : trapd;
  /* TG68KdotC_Kernel.vhd:3257:25  */
  assign n8006_o = clkena_lw ? next_micro_state : micro_state;
  /* TG68KdotC_Kernel.vhd:3255:17  */
  assign n8007_o = reset ? trapd : n8005_o;
  /* TG68KdotC_Kernel.vhd:3255:17  */
  assign n8009_o = reset ? 7'b0000010 : n8006_o;
  /* TG68KdotC_Kernel.vhd:3264:33  */
  assign n8015_o = micro_state == 7'b0000010;
  /* TG68KdotC_Kernel.vhd:3269:33  */
  assign n8018_o = micro_state == 7'b0000011;
  /* TG68KdotC_Kernel.vhd:3274:33  */
  assign n8021_o = micro_state == 7'b0000100;
  /* TG68KdotC_Kernel.vhd:3280:49  */
  assign n8022_o = brief[8];
  /* TG68KdotC_Kernel.vhd:3280:52  */
  assign n8023_o = ~n8022_o;
  /* TG68KdotC_Kernel.vhd:3280:57  */
  assign n8025_o = n8023_o | 1'b0;
  /* TG68KdotC_Kernel.vhd:3280:82  */
  assign n8026_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:3280:85  */
  assign n8027_o = ~n8026_o;
  /* TG68KdotC_Kernel.vhd:3280:90  */
  assign n8029_o = 1'b1 & n8027_o;
  /* TG68KdotC_Kernel.vhd:3280:75  */
  assign n8030_o = n8025_o | n8029_o;
  /* TG68KdotC_Kernel.vhd:3287:57  */
  assign n8032_o = brief[7];
  /* TG68KdotC_Kernel.vhd:3289:59  */
  assign n8033_o = exec[22];
  /* TG68KdotC_Kernel.vhd:3289:49  */
  assign n8035_o = n8033_o ? 1'b1 : n2164_o;
  /* TG68KdotC_Kernel.vhd:3287:49  */
  assign n8037_o = n8032_o ? 1'b1 : n2157_o;
  /* TG68KdotC_Kernel.vhd:3287:49  */
  assign n8038_o = n8032_o ? n2164_o : n8035_o;
  /* TG68KdotC_Kernel.vhd:3292:57  */
  assign n8039_o = brief[5];
  /* TG68KdotC_Kernel.vhd:3292:60  */
  assign n8040_o = ~n8039_o;
  /* TG68KdotC_Kernel.vhd:3295:65  */
  assign n8041_o = brief[4];
  assign n8043_o = n7810_o[0];
  assign n8044_o = n7782_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8045_o = n2184_o ? n8043_o : n8044_o;
  /* TG68KdotC_Kernel.vhd:3295:57  */
  assign n8046_o = n8041_o ? 1'b1 : n8045_o;
  /* TG68KdotC_Kernel.vhd:3292:49  */
  assign n8048_o = n8040_o ? 2'b01 : n7921_o;
  assign n8049_o = n7810_o[0];
  assign n8050_o = n7782_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8051_o = n2184_o ? n8049_o : n8050_o;
  /* TG68KdotC_Kernel.vhd:3292:49  */
  assign n8052_o = n8040_o ? n8051_o : n8046_o;
  /* TG68KdotC_Kernel.vhd:3280:41  */
  assign n8054_o = n8030_o ? 2'b01 : n8048_o;
  /* TG68KdotC_Kernel.vhd:3280:41  */
  assign n8057_o = n8030_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3280:41  */
  assign n8060_o = n8030_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3280:41  */
  assign n8061_o = n8030_o ? n2157_o : n8037_o;
  /* TG68KdotC_Kernel.vhd:3280:41  */
  assign n8062_o = n8030_o ? n2164_o : n8038_o;
  /* TG68KdotC_Kernel.vhd:3280:41  */
  assign n8063_o = n8030_o ? 1'b1 : n7832_o;
  assign n8064_o = n7810_o[0];
  assign n8065_o = n7782_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8066_o = n2184_o ? n8064_o : n8065_o;
  /* TG68KdotC_Kernel.vhd:3280:41  */
  assign n8067_o = n8030_o ? n8066_o : n8052_o;
  /* TG68KdotC_Kernel.vhd:3280:41  */
  assign n8070_o = n8030_o ? 7'b0000110 : 7'b0001011;
  /* TG68KdotC_Kernel.vhd:3279:33  */
  assign n8072_o = micro_state == 7'b0000101;
  /* TG68KdotC_Kernel.vhd:3302:33  */
  assign n8075_o = micro_state == 7'b0000110;
  /* TG68KdotC_Kernel.vhd:3310:49  */
  assign n8076_o = brief[5];
  /* TG68KdotC_Kernel.vhd:3310:41  */
  assign n8079_o = n8076_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3313:49  */
  assign n8080_o = brief[6];
  /* TG68KdotC_Kernel.vhd:3313:52  */
  assign n8081_o = ~n8080_o;
  /* TG68KdotC_Kernel.vhd:3313:66  */
  assign n8082_o = brief[2];
  /* TG68KdotC_Kernel.vhd:3313:69  */
  assign n8083_o = ~n8082_o;
  /* TG68KdotC_Kernel.vhd:3313:57  */
  assign n8084_o = n8083_o & n8081_o;
  /* TG68KdotC_Kernel.vhd:3316:57  */
  assign n8086_o = brief[1:0];
  /* TG68KdotC_Kernel.vhd:3316:69  */
  assign n8088_o = n8086_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:3316:49  */
  assign n8091_o = n8088_o ? 7'b0000110 : 7'b0001100;
  /* TG68KdotC_Kernel.vhd:3322:57  */
  assign n8092_o = brief[1:0];
  /* TG68KdotC_Kernel.vhd:3322:69  */
  assign n8094_o = n8092_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:3322:49  */
  assign n8098_o = n8094_o ? n7921_o : 2'b10;
  /* TG68KdotC_Kernel.vhd:3322:49  */
  assign n8101_o = n8094_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3322:49  */
  assign n8103_o = n8094_o ? 1'b1 : n7690_o;
  /* TG68KdotC_Kernel.vhd:3322:49  */
  assign n8104_o = n8094_o ? 1'b1 : n2170_o;
  assign n8105_o = n7810_o[0];
  assign n8106_o = n7782_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8107_o = n2184_o ? n8105_o : n8106_o;
  /* TG68KdotC_Kernel.vhd:3322:49  */
  assign n8108_o = n8094_o ? n8107_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3322:49  */
  assign n8110_o = n8094_o ? n7937_o : 7'b0001101;
  /* TG68KdotC_Kernel.vhd:3313:41  */
  assign n8112_o = n8084_o ? 2'b01 : n8098_o;
  /* TG68KdotC_Kernel.vhd:3313:41  */
  assign n8114_o = n8084_o ? 1'b0 : n8101_o;
  /* TG68KdotC_Kernel.vhd:3313:41  */
  assign n8115_o = n8084_o ? n7690_o : n8103_o;
  /* TG68KdotC_Kernel.vhd:3313:41  */
  assign n8116_o = n8084_o ? n2170_o : n8104_o;
  /* TG68KdotC_Kernel.vhd:3313:41  */
  assign n8117_o = n8084_o ? 1'b1 : n7832_o;
  assign n8118_o = n7810_o[0];
  assign n8119_o = n7782_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8120_o = n2184_o ? n8118_o : n8119_o;
  /* TG68KdotC_Kernel.vhd:3313:41  */
  assign n8121_o = n8084_o ? n8120_o : n8108_o;
  /* TG68KdotC_Kernel.vhd:3313:41  */
  assign n8122_o = n8084_o ? n8091_o : n8110_o;
  /* TG68KdotC_Kernel.vhd:3309:33  */
  assign n8124_o = micro_state == 7'b0001011;
  /* TG68KdotC_Kernel.vhd:3333:33  */
  assign n8127_o = micro_state == 7'b0001100;
  /* TG68KdotC_Kernel.vhd:3343:49  */
  assign n8129_o = brief[1];
  /* TG68KdotC_Kernel.vhd:3343:52  */
  assign n8130_o = ~n8129_o;
  /* TG68KdotC_Kernel.vhd:3346:57  */
  assign n8131_o = brief[0];
  assign n8133_o = n7810_o[0];
  assign n8134_o = n7782_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8135_o = n2184_o ? n8133_o : n8134_o;
  /* TG68KdotC_Kernel.vhd:3346:49  */
  assign n8136_o = n8131_o ? 1'b1 : n8135_o;
  /* TG68KdotC_Kernel.vhd:3343:41  */
  assign n8138_o = n8130_o ? 2'b01 : n7921_o;
  assign n8139_o = n7810_o[0];
  assign n8140_o = n7782_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8141_o = n2184_o ? n8139_o : n8140_o;
  /* TG68KdotC_Kernel.vhd:3343:41  */
  assign n8142_o = n8130_o ? n8141_o : n8136_o;
  /* TG68KdotC_Kernel.vhd:3340:33  */
  assign n8144_o = micro_state == 7'b0001101;
  /* TG68KdotC_Kernel.vhd:3353:49  */
  assign n8145_o = brief[1];
  /* TG68KdotC_Kernel.vhd:3353:41  */
  assign n8148_o = n8145_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3356:49  */
  assign n8149_o = brief[6];
  /* TG68KdotC_Kernel.vhd:3356:52  */
  assign n8150_o = ~n8149_o;
  /* TG68KdotC_Kernel.vhd:3356:66  */
  assign n8151_o = brief[2];
  /* TG68KdotC_Kernel.vhd:3356:57  */
  assign n8152_o = n8151_o & n8150_o;
  /* TG68KdotC_Kernel.vhd:3356:41  */
  assign n8156_o = n8152_o ? 2'b01 : n7921_o;
  /* TG68KdotC_Kernel.vhd:3356:41  */
  assign n8158_o = n8152_o ? n7690_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3356:41  */
  assign n8159_o = n8152_o ? n2170_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3356:41  */
  assign n8160_o = n8152_o ? 1'b1 : n7832_o;
  /* TG68KdotC_Kernel.vhd:3356:41  */
  assign n8162_o = n8152_o ? 7'b0000110 : n7937_o;
  /* TG68KdotC_Kernel.vhd:3352:33  */
  assign n8164_o = micro_state == 7'b0001110;
  /* TG68KdotC_Kernel.vhd:3366:33  */
  assign n8166_o = micro_state == 7'b0000111;
  /* TG68KdotC_Kernel.vhd:3372:49  */
  assign n8167_o = brief[8];
  /* TG68KdotC_Kernel.vhd:3372:52  */
  assign n8168_o = ~n8167_o;
  /* TG68KdotC_Kernel.vhd:3372:57  */
  assign n8170_o = n8168_o | 1'b0;
  /* TG68KdotC_Kernel.vhd:3372:82  */
  assign n8171_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:3372:85  */
  assign n8172_o = ~n8171_o;
  /* TG68KdotC_Kernel.vhd:3372:90  */
  assign n8174_o = 1'b1 & n8172_o;
  /* TG68KdotC_Kernel.vhd:3372:75  */
  assign n8175_o = n8170_o | n8174_o;
  /* TG68KdotC_Kernel.vhd:3379:57  */
  assign n8177_o = brief[7];
  /* TG68KdotC_Kernel.vhd:3379:49  */
  assign n8179_o = n8177_o ? 1'b1 : n2157_o;
  /* TG68KdotC_Kernel.vhd:3384:57  */
  assign n8180_o = brief[5];
  /* TG68KdotC_Kernel.vhd:3384:60  */
  assign n8181_o = ~n8180_o;
  /* TG68KdotC_Kernel.vhd:3387:65  */
  assign n8182_o = brief[4];
  assign n8184_o = n7810_o[0];
  assign n8185_o = n7782_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8186_o = n2184_o ? n8184_o : n8185_o;
  /* TG68KdotC_Kernel.vhd:3387:57  */
  assign n8187_o = n8182_o ? 1'b1 : n8186_o;
  /* TG68KdotC_Kernel.vhd:3384:49  */
  assign n8189_o = n8181_o ? 2'b01 : n7921_o;
  assign n8190_o = n7810_o[0];
  assign n8191_o = n7782_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8192_o = n2184_o ? n8190_o : n8191_o;
  /* TG68KdotC_Kernel.vhd:3384:49  */
  assign n8193_o = n8181_o ? n8192_o : n8187_o;
  /* TG68KdotC_Kernel.vhd:3372:41  */
  assign n8195_o = n8175_o ? 2'b01 : n8189_o;
  /* TG68KdotC_Kernel.vhd:3372:41  */
  assign n8198_o = n8175_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3372:41  */
  assign n8201_o = n8175_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3372:41  */
  assign n8202_o = n8175_o ? n2157_o : n8179_o;
  /* TG68KdotC_Kernel.vhd:3372:41  */
  assign n8203_o = n8175_o ? 1'b1 : n7832_o;
  assign n8204_o = n7810_o[0];
  assign n8205_o = n7782_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8206_o = n2184_o ? n8204_o : n8205_o;
  /* TG68KdotC_Kernel.vhd:3372:41  */
  assign n8207_o = n8175_o ? n8206_o : n8193_o;
  /* TG68KdotC_Kernel.vhd:3372:41  */
  assign n8210_o = n8175_o ? 7'b0010100 : 7'b0001111;
  /* TG68KdotC_Kernel.vhd:3371:33  */
  assign n8212_o = micro_state == 7'b0010011;
  /* TG68KdotC_Kernel.vhd:3394:33  */
  assign n8215_o = micro_state == 7'b0010100;
  /* TG68KdotC_Kernel.vhd:3403:49  */
  assign n8216_o = brief[5];
  /* TG68KdotC_Kernel.vhd:3403:41  */
  assign n8219_o = n8216_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3406:49  */
  assign n8220_o = brief[6];
  /* TG68KdotC_Kernel.vhd:3406:52  */
  assign n8221_o = ~n8220_o;
  /* TG68KdotC_Kernel.vhd:3406:66  */
  assign n8222_o = brief[2];
  /* TG68KdotC_Kernel.vhd:3406:69  */
  assign n8223_o = ~n8222_o;
  /* TG68KdotC_Kernel.vhd:3406:57  */
  assign n8224_o = n8223_o & n8221_o;
  /* TG68KdotC_Kernel.vhd:3409:57  */
  assign n8226_o = brief[1:0];
  /* TG68KdotC_Kernel.vhd:3409:69  */
  assign n8228_o = n8226_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:3409:49  */
  assign n8231_o = n8228_o ? 7'b0010100 : 7'b0010000;
  /* TG68KdotC_Kernel.vhd:3415:57  */
  assign n8232_o = brief[1:0];
  /* TG68KdotC_Kernel.vhd:3415:69  */
  assign n8234_o = n8232_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:3415:49  */
  assign n8239_o = n8234_o ? 2'b11 : 2'b10;
  assign n8240_o = n7803_o[1];
  assign n8241_o = n7601_o[1];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8242_o = n2184_o ? n8240_o : n8241_o;
  /* TG68KdotC_Kernel.vhd:3415:49  */
  assign n8243_o = n8234_o ? n8242_o : 1'b1;
  assign n8244_o = n7810_o[0];
  assign n8245_o = n7782_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8246_o = n2184_o ? n8244_o : n8245_o;
  /* TG68KdotC_Kernel.vhd:3415:49  */
  assign n8247_o = n8234_o ? n8246_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3415:49  */
  assign n8250_o = n8234_o ? 7'b0000001 : 7'b0010001;
  /* TG68KdotC_Kernel.vhd:3406:41  */
  assign n8252_o = n8224_o ? 2'b01 : n8239_o;
  assign n8253_o = n7803_o[1];
  assign n8254_o = n7601_o[1];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8255_o = n2184_o ? n8253_o : n8254_o;
  /* TG68KdotC_Kernel.vhd:3406:41  */
  assign n8256_o = n8224_o ? n8255_o : n8243_o;
  /* TG68KdotC_Kernel.vhd:3406:41  */
  assign n8257_o = n8224_o ? 1'b1 : n7832_o;
  assign n8258_o = n7810_o[0];
  assign n8259_o = n7782_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8260_o = n2184_o ? n8258_o : n8259_o;
  /* TG68KdotC_Kernel.vhd:3406:41  */
  assign n8261_o = n8224_o ? n8260_o : n8247_o;
  /* TG68KdotC_Kernel.vhd:3406:41  */
  assign n8262_o = n8224_o ? n8231_o : n8250_o;
  /* TG68KdotC_Kernel.vhd:3402:33  */
  assign n8264_o = micro_state == 7'b0001111;
  /* TG68KdotC_Kernel.vhd:3426:33  */
  assign n8268_o = micro_state == 7'b0010000;
  /* TG68KdotC_Kernel.vhd:3437:49  */
  assign n8271_o = brief[1];
  /* TG68KdotC_Kernel.vhd:3437:52  */
  assign n8272_o = ~n8271_o;
  /* TG68KdotC_Kernel.vhd:3440:57  */
  assign n8273_o = brief[0];
  assign n8275_o = n7810_o[0];
  assign n8276_o = n7782_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8277_o = n2184_o ? n8275_o : n8276_o;
  /* TG68KdotC_Kernel.vhd:3440:49  */
  assign n8278_o = n8273_o ? 1'b1 : n8277_o;
  /* TG68KdotC_Kernel.vhd:3437:41  */
  assign n8280_o = n8272_o ? 2'b01 : n7921_o;
  assign n8281_o = n7810_o[0];
  assign n8282_o = n7782_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8283_o = n2184_o ? n8281_o : n8282_o;
  /* TG68KdotC_Kernel.vhd:3437:41  */
  assign n8284_o = n8272_o ? n8283_o : n8278_o;
  /* TG68KdotC_Kernel.vhd:3433:33  */
  assign n8286_o = micro_state == 7'b0010001;
  /* TG68KdotC_Kernel.vhd:3448:49  */
  assign n8288_o = brief[1];
  /* TG68KdotC_Kernel.vhd:3448:41  */
  assign n8291_o = n8288_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3451:49  */
  assign n8292_o = brief[6];
  /* TG68KdotC_Kernel.vhd:3451:52  */
  assign n8293_o = ~n8292_o;
  /* TG68KdotC_Kernel.vhd:3451:66  */
  assign n8294_o = brief[2];
  /* TG68KdotC_Kernel.vhd:3451:57  */
  assign n8295_o = n8294_o & n8293_o;
  /* TG68KdotC_Kernel.vhd:3451:41  */
  assign n8299_o = n8295_o ? 2'b01 : 2'b11;
  /* TG68KdotC_Kernel.vhd:3451:41  */
  assign n8300_o = n8295_o ? 1'b1 : n7832_o;
  /* TG68KdotC_Kernel.vhd:3451:41  */
  assign n8303_o = n8295_o ? 7'b0010100 : 7'b0000001;
  /* TG68KdotC_Kernel.vhd:3446:33  */
  assign n8305_o = micro_state == 7'b0010010;
  /* TG68KdotC_Kernel.vhd:3462:41  */
  assign n8307_o = exe_condition ? 1'b1 : n7686_o;
  /* TG68KdotC_Kernel.vhd:3462:41  */
  assign n8310_o = exe_condition ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3462:41  */
  assign n8312_o = exe_condition ? 7'b0000001 : n7937_o;
  /* TG68KdotC_Kernel.vhd:3461:33  */
  assign n8314_o = micro_state == 7'b0010101;
  /* TG68KdotC_Kernel.vhd:3468:33  */
  assign n8316_o = micro_state == 7'b0010110;
  /* TG68KdotC_Kernel.vhd:3473:54  */
  assign n8317_o = ~long_start;
  /* TG68KdotC_Kernel.vhd:3473:41  */
  assign n8320_o = n8317_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3472:33  */
  assign n8323_o = micro_state == 7'b0010111;
  /* TG68KdotC_Kernel.vhd:3482:33  */
  assign n8325_o = micro_state == 7'b0011000;
  /* TG68KdotC_Kernel.vhd:3486:57  */
  assign n8326_o = ~exe_condition;
  /* TG68KdotC_Kernel.vhd:3488:57  */
  assign n8327_o = c_out[1];
  /* TG68KdotC_Kernel.vhd:3486:41  */
  assign n8329_o = n8335_o ? 1'b1 : n7686_o;
  /* TG68KdotC_Kernel.vhd:3488:49  */
  assign n8332_o = n8327_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3486:41  */
  assign n8334_o = n8341_o ? 7'b0000001 : n7937_o;
  /* TG68KdotC_Kernel.vhd:3486:41  */
  assign n8335_o = n8327_o & n8326_o;
  /* TG68KdotC_Kernel.vhd:3486:41  */
  assign n8338_o = n8326_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3486:41  */
  assign n8340_o = n8326_o ? n8332_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3486:41  */
  assign n8341_o = n8327_o & n8326_o;
  /* TG68KdotC_Kernel.vhd:3485:33  */
  assign n8343_o = micro_state == 7'b0011001;
  /* TG68KdotC_Kernel.vhd:3495:33  */
  assign n8349_o = micro_state == 7'b1001000;
  /* TG68KdotC_Kernel.vhd:3504:50  */
  assign n8350_o = sndopc[15];
  /* TG68KdotC_Kernel.vhd:3507:58  */
  assign n8351_o = opcode[10:9];
  /* TG68KdotC_Kernel.vhd:3507:71  */
  assign n8353_o = n8351_o == 2'b00;
  assign n8355_o = n1909_o[88];
  /* TG68KdotC_Kernel.vhd:3504:41  */
  assign n8356_o = n8363_o ? 1'b1 : n8355_o;
  /* TG68KdotC_Kernel.vhd:3504:41  */
  assign n8358_o = n8350_o ? 2'b10 : n7688_o;
  /* TG68KdotC_Kernel.vhd:3504:41  */
  assign n8361_o = n8350_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3504:41  */
  assign n8363_o = n8353_o & n8350_o;
  /* TG68KdotC_Kernel.vhd:3502:33  */
  assign n8368_o = micro_state == 7'b1001001;
  /* TG68KdotC_Kernel.vhd:3519:50  */
  assign n8370_o = sndopc[15];
  /* TG68KdotC_Kernel.vhd:3519:41  */
  assign n8372_o = n8370_o ? 2'b10 : n7688_o;
  /* TG68KdotC_Kernel.vhd:3519:41  */
  assign n8375_o = n8370_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3526:61  */
  assign n8379_o = exec[88];
  /* TG68KdotC_Kernel.vhd:3527:50  */
  assign n8380_o = sndopc[11];
  /* TG68KdotC_Kernel.vhd:3527:41  */
  assign n8382_o = n8380_o ? 2'b01 : n7921_o;
  /* TG68KdotC_Kernel.vhd:3527:41  */
  assign n8384_o = n8380_o ? 7'b1001011 : n7937_o;
  /* TG68KdotC_Kernel.vhd:3516:33  */
  assign n8386_o = micro_state == 7'b1001010;
  /* TG68KdotC_Kernel.vhd:3531:33  */
  assign n8388_o = micro_state == 7'b1001011;
  /* TG68KdotC_Kernel.vhd:3535:49  */
  assign n8389_o = flags[0];
  /* TG68KdotC_Kernel.vhd:3535:41  */
  assign n8391_o = n8389_o ? 1'b1 : n8003_o;
  /* TG68KdotC_Kernel.vhd:3534:33  */
  assign n8393_o = micro_state == 7'b1001100;
  /* TG68KdotC_Kernel.vhd:3540:33  */
  assign n8395_o = micro_state == 7'b0111110;
  /* TG68KdotC_Kernel.vhd:3545:49  */
  assign n8396_o = flags[2];
  /* TG68KdotC_Kernel.vhd:3545:41  */
  assign n8403_o = n8396_o ? 2'b11 : n7921_o;
  /* TG68KdotC_Kernel.vhd:3545:41  */
  assign n8406_o = n8396_o ? 1'b0 : 1'b1;
  assign n8407_o = n1909_o[27];
  /* TG68KdotC_Kernel.vhd:3545:41  */
  assign n8408_o = n8396_o ? n8407_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3545:41  */
  assign n8409_o = n8396_o ? n7795_o : 1'b1;
  assign n8410_o = n7797_o[4];
  assign n8411_o = n7779_o[4];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8412_o = n2184_o ? n8410_o : n8411_o;
  /* TG68KdotC_Kernel.vhd:3545:41  */
  assign n8413_o = n8396_o ? 1'b1 : n8412_o;
  /* TG68KdotC_Kernel.vhd:3545:41  */
  assign n8414_o = n8396_o ? 1'b1 : n1925_o;
  assign n8415_o = n1909_o[85];
  assign n8416_o = n7783_o[1];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8417_o = n2184_o ? n8415_o : n8416_o;
  /* TG68KdotC_Kernel.vhd:3545:41  */
  assign n8418_o = n8396_o ? n8417_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3545:41  */
  assign n8420_o = n8396_o ? 7'b0000001 : n7937_o;
  /* TG68KdotC_Kernel.vhd:3543:33  */
  assign n8422_o = micro_state == 7'b0111111;
  /* TG68KdotC_Kernel.vhd:3559:63  */
  assign n8423_o = sndopc[15];
  /* TG68KdotC_Kernel.vhd:3557:33  */
  assign n8426_o = micro_state == 7'b1000000;
  /* TG68KdotC_Kernel.vhd:3562:33  */
  assign n8432_o = micro_state == 7'b1000001;
  /* TG68KdotC_Kernel.vhd:3570:33  */
  assign n8435_o = micro_state == 7'b1000010;
  /* TG68KdotC_Kernel.vhd:3575:49  */
  assign n8436_o = flags[2];
  assign n8438_o = n1909_o[86];
  assign n8439_o = n7783_o[2];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8440_o = n2184_o ? n8438_o : n8439_o;
  /* TG68KdotC_Kernel.vhd:3575:41  */
  assign n8441_o = n8436_o ? 1'b1 : n8440_o;
  /* TG68KdotC_Kernel.vhd:3574:33  */
  assign n8447_o = micro_state == 7'b1000011;
  /* TG68KdotC_Kernel.vhd:3585:33  */
  assign n8450_o = micro_state == 7'b1000100;
  /* TG68KdotC_Kernel.vhd:3590:49  */
  assign n8451_o = flags[2];
  /* TG68KdotC_Kernel.vhd:3594:71  */
  assign n8453_o = sndopc[15];
  /* TG68KdotC_Kernel.vhd:3590:41  */
  assign n8461_o = n8451_o ? 2'b11 : n7921_o;
  /* TG68KdotC_Kernel.vhd:3590:41  */
  assign n8464_o = n8451_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3590:41  */
  assign n8466_o = n8451_o ? n8453_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:3590:41  */
  assign n8469_o = n8451_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:3590:41  */
  assign n8471_o = n8451_o ? 1'b1 : n7727_o;
  assign n8472_o = n1909_o[27];
  /* TG68KdotC_Kernel.vhd:3590:41  */
  assign n8473_o = n8451_o ? n8472_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3590:41  */
  assign n8474_o = n8451_o ? n7795_o : 1'b1;
  assign n8475_o = n7797_o[4];
  assign n8476_o = n7779_o[4];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8477_o = n2184_o ? n8475_o : n8476_o;
  /* TG68KdotC_Kernel.vhd:3590:41  */
  assign n8478_o = n8451_o ? 1'b1 : n8477_o;
  /* TG68KdotC_Kernel.vhd:3590:41  */
  assign n8479_o = n8451_o ? 1'b1 : n2170_o;
  assign n8480_o = n7803_o[1];
  assign n8481_o = n7601_o[1];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8482_o = n2184_o ? n8480_o : n8481_o;
  /* TG68KdotC_Kernel.vhd:3590:41  */
  assign n8483_o = n8451_o ? n8482_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3590:41  */
  assign n8484_o = n8451_o ? n7815_o : 1'b1;
  assign n8485_o = n1909_o[85];
  assign n8486_o = n7783_o[1];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8487_o = n2184_o ? n8485_o : n8486_o;
  /* TG68KdotC_Kernel.vhd:3590:41  */
  assign n8488_o = n8451_o ? n8487_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3590:41  */
  assign n8491_o = n8451_o ? 7'b1000110 : 7'b1000111;
  /* TG68KdotC_Kernel.vhd:3589:33  */
  assign n8493_o = micro_state == 7'b1000101;
  /* TG68KdotC_Kernel.vhd:3607:33  */
  assign n8497_o = micro_state == 7'b1000110;
  /* TG68KdotC_Kernel.vhd:3614:33  */
  assign n8501_o = micro_state == 7'b1000111;
  /* TG68KdotC_Kernel.vhd:3620:58  */
  assign n8502_o = last_data_read[15:0];
  /* TG68KdotC_Kernel.vhd:3620:71  */
  assign n8504_o = n8502_o != 16'b0000000000000000;
  /* TG68KdotC_Kernel.vhd:3622:58  */
  assign n8505_o = opcode[5:3];
  /* TG68KdotC_Kernel.vhd:3622:70  */
  assign n8507_o = n8505_o == 3'b100;
  /* TG68KdotC_Kernel.vhd:3624:63  */
  assign n8509_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:3620:41  */
  assign n8511_o = n8519_o ? 1'b1 : n7795_o;
  /* TG68KdotC_Kernel.vhd:3622:49  */
  assign n8512_o = n8509_o & n8507_o;
  assign n8513_o = n7801_o[9];
  assign n8514_o = n7781_o[9];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8515_o = n2184_o ? n8513_o : n8514_o;
  /* TG68KdotC_Kernel.vhd:3622:49  */
  assign n8516_o = n8507_o ? 1'b1 : n8515_o;
  /* TG68KdotC_Kernel.vhd:3620:41  */
  assign n8518_o = n8504_o ? 2'b01 : n7921_o;
  /* TG68KdotC_Kernel.vhd:3620:41  */
  assign n8519_o = n8512_o & n8504_o;
  assign n8520_o = n7801_o[9];
  assign n8521_o = n7781_o[9];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8522_o = n2184_o ? n8520_o : n8521_o;
  /* TG68KdotC_Kernel.vhd:3620:41  */
  assign n8523_o = n8504_o ? n8516_o : n8522_o;
  /* TG68KdotC_Kernel.vhd:3620:41  */
  assign n8525_o = n8504_o ? 7'b0011011 : n7937_o;
  /* TG68KdotC_Kernel.vhd:3619:33  */
  assign n8527_o = micro_state == 7'b0011010;
  /* TG68KdotC_Kernel.vhd:3631:53  */
  assign n8528_o = ~movem_run;
  /* TG68KdotC_Kernel.vhd:3637:58  */
  assign n8531_o = opcode[10];
  /* TG68KdotC_Kernel.vhd:3637:62  */
  assign n8532_o = ~n8531_o;
  /* TG68KdotC_Kernel.vhd:3637:49  */
  assign n8536_o = n8532_o ? 2'b11 : 2'b10;
  assign n8537_o = n7797_o[4];
  assign n8538_o = n7779_o[4];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8539_o = n2184_o ? n8537_o : n8538_o;
  /* TG68KdotC_Kernel.vhd:3637:49  */
  assign n8540_o = n8532_o ? 1'b1 : n8539_o;
  /* TG68KdotC_Kernel.vhd:3631:41  */
  assign n8542_o = n8528_o ? 2'b01 : n8536_o;
  assign n8543_o = n7797_o[4];
  assign n8544_o = n7779_o[4];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8545_o = n2184_o ? n8543_o : n8544_o;
  /* TG68KdotC_Kernel.vhd:3631:41  */
  assign n8546_o = n8528_o ? n8545_o : n8540_o;
  assign n8547_o = n7801_o[9];
  assign n8548_o = n7781_o[9];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8549_o = n2184_o ? n8547_o : n8548_o;
  /* TG68KdotC_Kernel.vhd:3631:41  */
  assign n8550_o = n8528_o ? n8549_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3631:41  */
  assign n8551_o = n8528_o ? n7806_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3631:41  */
  assign n8553_o = n8528_o ? n7937_o : 7'b0011011;
  /* TG68KdotC_Kernel.vhd:3630:33  */
  assign n8555_o = micro_state == 7'b0011011;
  /* TG68KdotC_Kernel.vhd:3646:50  */
  assign n8556_o = opcode[5:4];
  /* TG68KdotC_Kernel.vhd:3646:62  */
  assign n8558_o = n8556_o != 2'b00;
  /* TG68KdotC_Kernel.vhd:3646:41  */
  assign n8560_o = n8558_o ? 1'b1 : n7690_o;
  /* TG68KdotC_Kernel.vhd:3645:33  */
  assign n8562_o = micro_state == 7'b0011101;
  /* TG68KdotC_Kernel.vhd:3651:50  */
  assign n8563_o = opcode[2:0];
  /* TG68KdotC_Kernel.vhd:3651:62  */
  assign n8565_o = n8563_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:3651:41  */
  assign n8567_o = n8565_o ? 1'b1 : n7975_o;
  /* TG68KdotC_Kernel.vhd:3650:33  */
  assign n8572_o = micro_state == 7'b0011110;
  /* TG68KdotC_Kernel.vhd:3661:50  */
  assign n8573_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:3661:63  */
  assign n8575_o = n8573_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:3661:41  */
  assign n8577_o = n8575_o ? 1'b1 : n7975_o;
  /* TG68KdotC_Kernel.vhd:3666:50  */
  assign n8579_o = opcode[7:6];
  /* TG68KdotC_Kernel.vhd:3666:63  */
  assign n8581_o = n8579_o == 2'b01;
  /* TG68KdotC_Kernel.vhd:3666:41  */
  assign n8584_o = n8581_o ? 2'b00 : 2'b01;
  /* TG68KdotC_Kernel.vhd:3660:33  */
  assign n8587_o = micro_state == 7'b0011111;
  /* TG68KdotC_Kernel.vhd:3676:33  */
  assign n8589_o = micro_state == 7'b0100000;
  /* TG68KdotC_Kernel.vhd:3680:50  */
  assign n8590_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:3680:63  */
  assign n8592_o = n8590_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:3680:41  */
  assign n8594_o = n8592_o ? 1'b1 : n7975_o;
  /* TG68KdotC_Kernel.vhd:3679:33  */
  assign n8597_o = micro_state == 7'b0100001;
  /* TG68KdotC_Kernel.vhd:3690:50  */
  assign n8598_o = opcode[11:9];
  /* TG68KdotC_Kernel.vhd:3690:63  */
  assign n8600_o = n8598_o == 3'b111;
  /* TG68KdotC_Kernel.vhd:3690:41  */
  assign n8602_o = n8600_o ? 1'b1 : n7975_o;
  /* TG68KdotC_Kernel.vhd:3689:33  */
  assign n8605_o = micro_state == 7'b0100010;
  /* TG68KdotC_Kernel.vhd:3699:33  */
  assign n8609_o = micro_state == 7'b0100011;
  /* TG68KdotC_Kernel.vhd:3705:33  */
  assign n8612_o = micro_state == 7'b0100100;
  /* TG68KdotC_Kernel.vhd:3709:33  */
  assign n8615_o = micro_state == 7'b0100101;
  /* TG68KdotC_Kernel.vhd:3714:33  */
  assign n8618_o = micro_state == 7'b0100110;
  /* TG68KdotC_Kernel.vhd:3718:33  */
  assign n8621_o = micro_state == 7'b0110010;
  /* TG68KdotC_Kernel.vhd:3735:71  */
  assign n8624_o = trap_interrupt | trap_trace;
  /* TG68KdotC_Kernel.vhd:3735:89  */
  assign n8625_o = n8624_o | trap_berr;
  /* TG68KdotC_Kernel.vhd:3735:49  */
  assign n8627_o = n8625_o ? 1'b1 : n8000_o;
  /* TG68KdotC_Kernel.vhd:3729:41  */
  assign n8630_o = use_vbr_stackframe ? 2'b01 : 2'b10;
  /* TG68KdotC_Kernel.vhd:3729:41  */
  assign n8631_o = use_vbr_stackframe ? n8000_o : n8627_o;
  /* TG68KdotC_Kernel.vhd:3729:41  */
  assign n8632_o = use_vbr_stackframe ? 1'b1 : n1960_o;
  /* TG68KdotC_Kernel.vhd:3729:41  */
  assign n8635_o = use_vbr_stackframe ? 7'b0110100 : 7'b0110101;
  /* TG68KdotC_Kernel.vhd:3725:33  */
  assign n8637_o = micro_state == 7'b0110011;
  /* TG68KdotC_Kernel.vhd:3743:63  */
  assign n8638_o = trap_interrupt | trap_trace;
  /* TG68KdotC_Kernel.vhd:3743:41  */
  assign n8640_o = n8638_o ? 1'b1 : n8000_o;
  /* TG68KdotC_Kernel.vhd:3742:33  */
  assign n8643_o = micro_state == 7'b0110100;
  /* TG68KdotC_Kernel.vhd:3751:33  */
  assign n8646_o = micro_state == 7'b0110101;
  /* TG68KdotC_Kernel.vhd:3758:33  */
  assign n8650_o = micro_state == 7'b0110110;
  /* TG68KdotC_Kernel.vhd:3770:33  */
  assign n8653_o = micro_state == 7'b0110111;
  /* TG68KdotC_Kernel.vhd:3776:33  */
  assign n8656_o = micro_state == 7'b0111000;
  /* TG68KdotC_Kernel.vhd:3782:33  */
  assign n8659_o = micro_state == 7'b0111001;
  /* TG68KdotC_Kernel.vhd:3788:33  */
  assign n8662_o = micro_state == 7'b0111010;
  /* TG68KdotC_Kernel.vhd:3794:33  */
  assign n8665_o = micro_state == 7'b0111011;
  /* TG68KdotC_Kernel.vhd:3800:33  */
  assign n8668_o = micro_state == 7'b0111100;
  /* TG68KdotC_Kernel.vhd:3806:33  */
  assign n8671_o = micro_state == 7'b0111101;
  /* TG68KdotC_Kernel.vhd:3826:62  */
  assign n8674_o = ~use_vbr_stackframe;
  /* TG68KdotC_Kernel.vhd:3826:76  */
  assign n8675_o = opcode[2];
  /* TG68KdotC_Kernel.vhd:3826:67  */
  assign n8676_o = n8674_o | n8675_o;
  /* TG68KdotC_Kernel.vhd:3826:41  */
  assign n8679_o = n8676_o ? 1'b1 : n7827_o;
  assign n8680_o = n7801_o[12];
  assign n8681_o = n7781_o[12];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8682_o = n2184_o ? n8680_o : n8681_o;
  /* TG68KdotC_Kernel.vhd:3826:41  */
  assign n8683_o = n8676_o ? 1'b1 : n8682_o;
  /* TG68KdotC_Kernel.vhd:3820:33  */
  assign n8685_o = micro_state == 7'b0101011;
  /* TG68KdotC_Kernel.vhd:3834:77  */
  assign n8687_o = opcode[2];
  /* TG68KdotC_Kernel.vhd:3834:80  */
  assign n8688_o = ~n8687_o;
  /* TG68KdotC_Kernel.vhd:3834:67  */
  assign n8689_o = n8688_o & use_vbr_stackframe;
  /* TG68KdotC_Kernel.vhd:3834:41  */
  assign n8692_o = n8689_o ? 2'b10 : n7921_o;
  /* TG68KdotC_Kernel.vhd:3834:41  */
  assign n8694_o = n8689_o ? 1'b1 : n7701_o;
  /* TG68KdotC_Kernel.vhd:3834:41  */
  assign n8695_o = n8689_o ? 1'b1 : n7987_o;
  /* TG68KdotC_Kernel.vhd:3834:41  */
  assign n8698_o = n8689_o ? 7'b0101101 : 7'b0000001;
  /* TG68KdotC_Kernel.vhd:3831:33  */
  assign n8700_o = micro_state == 7'b0101100;
  /* TG68KdotC_Kernel.vhd:3847:33  */
  assign n8702_o = micro_state == 7'b0101101;
  /* TG68KdotC_Kernel.vhd:3854:56  */
  assign n8703_o = last_data_in[15:12];
  /* TG68KdotC_Kernel.vhd:3854:70  */
  assign n8705_o = n8703_o == 4'b0010;
  /* TG68KdotC_Kernel.vhd:3854:41  */
  assign n8709_o = n8705_o ? 2'b10 : 2'b01;
  /* TG68KdotC_Kernel.vhd:3854:41  */
  assign n8711_o = n8705_o ? 2'b10 : n7921_o;
  /* TG68KdotC_Kernel.vhd:3854:41  */
  assign n8713_o = n8705_o ? 1'b1 : n7701_o;
  /* TG68KdotC_Kernel.vhd:3854:41  */
  assign n8714_o = n8705_o ? 1'b1 : n7987_o;
  /* TG68KdotC_Kernel.vhd:3854:41  */
  assign n8717_o = n8705_o ? 7'b0101111 : 7'b0000001;
  /* TG68KdotC_Kernel.vhd:3852:33  */
  assign n8719_o = micro_state == 7'b0101110;
  /* TG68KdotC_Kernel.vhd:3865:33  */
  assign n8721_o = micro_state == 7'b0101111;
  /* TG68KdotC_Kernel.vhd:3869:33  */
  assign n8723_o = micro_state == 7'b0110000;
  /* TG68KdotC_Kernel.vhd:3871:33  */
  assign n8726_o = micro_state == 7'b0110001;
  /* TG68KdotC_Kernel.vhd:3878:50  */
  assign n8728_o = brief[11:0];
  /* TG68KdotC_Kernel.vhd:3878:63  */
  assign n8730_o = n8728_o == 12'b000000000000;
  /* TG68KdotC_Kernel.vhd:3878:79  */
  assign n8731_o = brief[11:0];
  /* TG68KdotC_Kernel.vhd:3878:92  */
  assign n8733_o = n8731_o == 12'b000000000001;
  /* TG68KdotC_Kernel.vhd:3878:71  */
  assign n8734_o = n8730_o | n8733_o;
  /* TG68KdotC_Kernel.vhd:3878:108  */
  assign n8735_o = brief[11:0];
  /* TG68KdotC_Kernel.vhd:3878:121  */
  assign n8737_o = n8735_o == 12'b100000000000;
  /* TG68KdotC_Kernel.vhd:3878:100  */
  assign n8738_o = n8734_o | n8737_o;
  /* TG68KdotC_Kernel.vhd:3878:137  */
  assign n8739_o = brief[11:0];
  /* TG68KdotC_Kernel.vhd:3878:150  */
  assign n8741_o = n8739_o == 12'b100000000001;
  /* TG68KdotC_Kernel.vhd:3878:129  */
  assign n8742_o = n8738_o | n8741_o;
  /* TG68KdotC_Kernel.vhd:3879:48  */
  assign n8743_o = cpu[1];
  /* TG68KdotC_Kernel.vhd:3879:66  */
  assign n8744_o = brief[11:0];
  /* TG68KdotC_Kernel.vhd:3879:79  */
  assign n8746_o = n8744_o == 12'b000000000010;
  /* TG68KdotC_Kernel.vhd:3879:95  */
  assign n8747_o = brief[11:0];
  /* TG68KdotC_Kernel.vhd:3879:108  */
  assign n8749_o = n8747_o == 12'b100000000010;
  /* TG68KdotC_Kernel.vhd:3879:87  */
  assign n8750_o = n8746_o | n8749_o;
  /* TG68KdotC_Kernel.vhd:3879:124  */
  assign n8751_o = brief[11:0];
  /* TG68KdotC_Kernel.vhd:3879:137  */
  assign n8753_o = n8751_o == 12'b100000000011;
  /* TG68KdotC_Kernel.vhd:3879:116  */
  assign n8754_o = n8750_o | n8753_o;
  /* TG68KdotC_Kernel.vhd:3879:153  */
  assign n8755_o = brief[11:0];
  /* TG68KdotC_Kernel.vhd:3879:166  */
  assign n8757_o = n8755_o == 12'b100000000100;
  /* TG68KdotC_Kernel.vhd:3879:145  */
  assign n8758_o = n8754_o | n8757_o;
  /* TG68KdotC_Kernel.vhd:3879:56  */
  assign n8759_o = n8758_o & n8743_o;
  /* TG68KdotC_Kernel.vhd:3878:159  */
  assign n8760_o = n8742_o | n8759_o;
  /* TG68KdotC_Kernel.vhd:3880:58  */
  assign n8761_o = opcode[0];
  /* TG68KdotC_Kernel.vhd:3880:61  */
  assign n8762_o = ~n8761_o;
  /* TG68KdotC_Kernel.vhd:3878:41  */
  assign n8764_o = n8769_o ? 1'b1 : n7795_o;
  /* TG68KdotC_Kernel.vhd:3878:41  */
  assign n8766_o = n8760_o ? n7740_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3878:41  */
  assign n8768_o = n8760_o ? n8003_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:3878:41  */
  assign n8769_o = n8762_o & n8760_o;
  /* TG68KdotC_Kernel.vhd:3875:33  */
  assign n8771_o = micro_state == 7'b1001101;
  /* TG68KdotC_Kernel.vhd:3896:50  */
  assign n8775_o = opcode[6];
  assign n8777_o = n7797_o[1];
  assign n8778_o = n7779_o[1];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8779_o = n2184_o ? n8777_o : n8778_o;
  /* TG68KdotC_Kernel.vhd:3896:41  */
  assign n8780_o = n8775_o ? 1'b1 : n8779_o;
  /* TG68KdotC_Kernel.vhd:3899:50  */
  assign n8781_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:3899:53  */
  assign n8782_o = ~n8781_o;
  /* TG68KdotC_Kernel.vhd:3899:41  */
  assign n8785_o = n8782_o ? 2'b10 : 2'b11;
  /* TG68KdotC_Kernel.vhd:3891:33  */
  assign n8787_o = micro_state == 7'b1001110;
  /* TG68KdotC_Kernel.vhd:3906:50  */
  assign n8788_o = opcode[6];
  assign n8791_o = n7797_o[3];
  assign n8792_o = n7779_o[3];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8793_o = n2184_o ? n8791_o : n8792_o;
  /* TG68KdotC_Kernel.vhd:3906:41  */
  assign n8794_o = n8788_o ? 1'b1 : n8793_o;
  assign n8795_o = n7801_o[9];
  assign n8796_o = n7781_o[9];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8797_o = n2184_o ? n8795_o : n8796_o;
  /* TG68KdotC_Kernel.vhd:3906:41  */
  assign n8798_o = n8788_o ? 1'b1 : n8797_o;
  /* TG68KdotC_Kernel.vhd:3910:50  */
  assign n8799_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:3910:53  */
  assign n8800_o = ~n8799_o;
  /* TG68KdotC_Kernel.vhd:3910:41  */
  assign n8803_o = n8800_o ? 2'b10 : 2'b11;
  /* TG68KdotC_Kernel.vhd:3905:33  */
  assign n8805_o = micro_state == 7'b1001111;
  /* TG68KdotC_Kernel.vhd:3917:50  */
  assign n8806_o = opcode[6];
  /* TG68KdotC_Kernel.vhd:3921:58  */
  assign n8810_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:3921:61  */
  assign n8811_o = ~n8810_o;
  /* TG68KdotC_Kernel.vhd:3921:49  */
  assign n8814_o = n8811_o ? 2'b10 : 2'b11;
  /* TG68KdotC_Kernel.vhd:3917:41  */
  assign n8816_o = n8806_o ? n7687_o : 2'b01;
  /* TG68KdotC_Kernel.vhd:3917:41  */
  assign n8817_o = n8806_o ? n8814_o : n7921_o;
  assign n8818_o = n7797_o[3];
  assign n8819_o = n7779_o[3];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8820_o = n2184_o ? n8818_o : n8819_o;
  /* TG68KdotC_Kernel.vhd:3917:41  */
  assign n8821_o = n8806_o ? 1'b1 : n8820_o;
  assign n8822_o = n7801_o[9];
  assign n8823_o = n7781_o[9];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8824_o = n2184_o ? n8822_o : n8823_o;
  /* TG68KdotC_Kernel.vhd:3917:41  */
  assign n8825_o = n8806_o ? 1'b1 : n8824_o;
  /* TG68KdotC_Kernel.vhd:3917:41  */
  assign n8826_o = n8806_o ? 1'b1 : n7831_o;
  /* TG68KdotC_Kernel.vhd:3917:41  */
  assign n8828_o = n8806_o ? 7'b1010001 : n7937_o;
  /* TG68KdotC_Kernel.vhd:3916:33  */
  assign n8830_o = micro_state == 7'b1010000;
  /* TG68KdotC_Kernel.vhd:3931:50  */
  assign n8831_o = opcode[7];
  /* TG68KdotC_Kernel.vhd:3931:53  */
  assign n8832_o = ~n8831_o;
  /* TG68KdotC_Kernel.vhd:3931:41  */
  assign n8835_o = n8832_o ? 2'b10 : 2'b11;
  /* TG68KdotC_Kernel.vhd:3930:33  */
  assign n8837_o = micro_state == 7'b1010001;
  /* TG68KdotC_Kernel.vhd:3937:33  */
  assign n8839_o = micro_state == 7'b1010010;
  /* TG68KdotC_Kernel.vhd:3941:50  */
  assign n8840_o = opcode[15];
  /* TG68KdotC_Kernel.vhd:3941:59  */
  assign n8842_o = n8840_o | 1'b0;
  /* TG68KdotC_Kernel.vhd:3941:41  */
  assign n8845_o = n8842_o ? 6'b001110 : 6'b011110;
  /* TG68KdotC_Kernel.vhd:3940:33  */
  assign n8847_o = micro_state == 7'b1010101;
  /* TG68KdotC_Kernel.vhd:3950:51  */
  assign n8850_o = rot_cnt == 6'b000001;
  /* TG68KdotC_Kernel.vhd:3950:41  */
  assign n8853_o = n8850_o ? 7'b1010111 : 7'b1010110;
  /* TG68KdotC_Kernel.vhd:3948:33  */
  assign n8855_o = micro_state == 7'b1010110;
  /* TG68KdotC_Kernel.vhd:3957:50  */
  assign n8856_o = opcode[15];
  /* TG68KdotC_Kernel.vhd:3957:54  */
  assign n8857_o = ~n8856_o;
  /* TG68KdotC_Kernel.vhd:3957:41  */
  assign n8859_o = n8857_o ? 1'b1 : n7815_o;
  /* TG68KdotC_Kernel.vhd:3962:50  */
  assign n8861_o = opcode[15];
  /* TG68KdotC_Kernel.vhd:3962:54  */
  assign n8862_o = ~n8861_o;
  /* TG68KdotC_Kernel.vhd:3962:59  */
  assign n8864_o = 1'b1 & n8862_o;
  /* TG68KdotC_Kernel.vhd:3965:58  */
  assign n8866_o = sndopc[10];
  /* TG68KdotC_Kernel.vhd:3962:41  */
  assign n8868_o = n8872_o ? 2'b01 : n7921_o;
  /* TG68KdotC_Kernel.vhd:3962:41  */
  assign n8870_o = n8878_o ? 7'b1011000 : n7937_o;
  /* TG68KdotC_Kernel.vhd:3962:41  */
  assign n8872_o = n8866_o & n8864_o;
  /* TG68KdotC_Kernel.vhd:3962:41  */
  assign n8874_o = n8864_o ? 1'b1 : n7727_o;
  /* TG68KdotC_Kernel.vhd:3962:41  */
  assign n8875_o = n8864_o ? 1'b1 : n7795_o;
  assign n8876_o = n1909_o[67];
  /* TG68KdotC_Kernel.vhd:3962:41  */
  assign n8877_o = n8864_o ? 1'b1 : n8876_o;
  /* TG68KdotC_Kernel.vhd:3962:41  */
  assign n8878_o = n8866_o & n8864_o;
  /* TG68KdotC_Kernel.vhd:3956:33  */
  assign n8880_o = micro_state == 7'b1010111;
  /* TG68KdotC_Kernel.vhd:3972:33  */
  assign n8885_o = micro_state == 7'b1011000;
  /* TG68KdotC_Kernel.vhd:3978:33  */
  assign n8887_o = micro_state == 7'b1011001;
  /* TG68KdotC_Kernel.vhd:3982:51  */
  assign n8888_o = op2out[31:16];
  /* TG68KdotC_Kernel.vhd:3982:65  */
  assign n8890_o = n8888_o == 16'b0000000000000000;
  /* TG68KdotC_Kernel.vhd:3982:83  */
  assign n8891_o = opcode[15];
  /* TG68KdotC_Kernel.vhd:3982:74  */
  assign n8892_o = n8890_o | n8891_o;
  /* TG68KdotC_Kernel.vhd:3982:92  */
  assign n8894_o = n8892_o | 1'b0;
  /* TG68KdotC_Kernel.vhd:3982:117  */
  assign n8895_o = op2out[15:0];
  /* TG68KdotC_Kernel.vhd:3982:130  */
  assign n8897_o = n8895_o == 16'b0000000000000000;
  /* TG68KdotC_Kernel.vhd:3982:107  */
  assign n8898_o = n8897_o & n8894_o;
  /* TG68KdotC_Kernel.vhd:3982:41  */
  assign n8901_o = n8898_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:3982:41  */
  assign n8903_o = n8898_o ? n7937_o : 7'b1011011;
  /* TG68KdotC_Kernel.vhd:3981:33  */
  assign n8906_o = micro_state == 7'b1011010;
  /* TG68KdotC_Kernel.vhd:3990:50  */
  assign n8907_o = opcode[15];
  /* TG68KdotC_Kernel.vhd:3990:59  */
  assign n8909_o = n8907_o | 1'b0;
  /* TG68KdotC_Kernel.vhd:3990:41  */
  assign n8912_o = n8909_o ? 6'b001101 : 6'b011101;
  /* TG68KdotC_Kernel.vhd:3989:33  */
  assign n8914_o = micro_state == 7'b1011011;
  /* TG68KdotC_Kernel.vhd:3999:51  */
  assign n8917_o = rot_cnt == 6'b000001;
  /* TG68KdotC_Kernel.vhd:3999:41  */
  assign n8920_o = n8917_o ? 7'b1011101 : 7'b1011100;
  /* TG68KdotC_Kernel.vhd:3997:33  */
  assign n8922_o = micro_state == 7'b1011100;
  /* TG68KdotC_Kernel.vhd:4005:51  */
  assign n8923_o = ~z_error;
  /* TG68KdotC_Kernel.vhd:4005:70  */
  assign n8924_o = ~set_v_flag;
  /* TG68KdotC_Kernel.vhd:4005:56  */
  assign n8925_o = n8924_o & n8923_o;
  /* TG68KdotC_Kernel.vhd:4005:41  */
  assign n8927_o = n8925_o ? 1'b1 : n7795_o;
  /* TG68KdotC_Kernel.vhd:4008:50  */
  assign n8928_o = opcode[15];
  /* TG68KdotC_Kernel.vhd:4008:54  */
  assign n8929_o = ~n8928_o;
  /* TG68KdotC_Kernel.vhd:4008:59  */
  assign n8931_o = 1'b1 & n8929_o;
  /* TG68KdotC_Kernel.vhd:4008:41  */
  assign n8934_o = n8931_o ? 2'b01 : n7921_o;
  /* TG68KdotC_Kernel.vhd:4008:41  */
  assign n8937_o = n8931_o ? 1'b1 : 1'b0;
  assign n8938_o = n1909_o[68];
  /* TG68KdotC_Kernel.vhd:4008:41  */
  assign n8939_o = n8931_o ? 1'b1 : n8938_o;
  /* TG68KdotC_Kernel.vhd:4008:41  */
  assign n8941_o = n8931_o ? 7'b1011110 : n7937_o;
  /* TG68KdotC_Kernel.vhd:4004:33  */
  assign n8944_o = micro_state == 7'b1011101;
  /* TG68KdotC_Kernel.vhd:4017:48  */
  assign n8945_o = exec[34];
  /* TG68KdotC_Kernel.vhd:4017:41  */
  assign n8948_o = n8945_o ? 1'b1 : n7795_o;
  assign n8949_o = n7801_o[3];
  assign n8950_o = n7781_o[3];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n8951_o = n2184_o ? n8949_o : n8950_o;
  /* TG68KdotC_Kernel.vhd:4017:41  */
  assign n8952_o = n8945_o ? n8951_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:4016:33  */
  assign n8955_o = micro_state == 7'b1011110;
  /* TG68KdotC_Kernel.vhd:4026:50  */
  assign n8956_o = op2out[5:0];
  /* TG68KdotC_Kernel.vhd:4026:62  */
  assign n8958_o = n8956_o != 6'b000000;
  /* TG68KdotC_Kernel.vhd:4027:70  */
  assign n8959_o = op2out[5:0];
  /* TG68KdotC_Kernel.vhd:4026:41  */
  assign n8961_o = n8958_o ? n8959_o : n7734_o;
  assign n8962_o = n7853_o[23];
  /* TG68KdotC_Kernel.vhd:4026:41  */
  assign n8963_o = n8958_o ? n8962_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:4025:33  */
  assign n8965_o = micro_state == 7'b1010011;
  /* TG68KdotC_Kernel.vhd:4032:33  */
  assign n8967_o = micro_state == 7'b1010100;
  assign n8968_o = {n8967_o, n8965_o, n8955_o, n8944_o, n8922_o, n8914_o, n8906_o, n8887_o, n8885_o, n8880_o, n8855_o, n8847_o, n8839_o, n8837_o, n8830_o, n8805_o, n8787_o, n8771_o, n8726_o, n8723_o, n8721_o, n8719_o, n8702_o, n8700_o, n8685_o, n8671_o, n8668_o, n8665_o, n8662_o, n8659_o, n8656_o, n8653_o, n8650_o, n8646_o, n8643_o, n8637_o, n8621_o, n8618_o, n8615_o, n8612_o, n8609_o, n8605_o, n8597_o, n8589_o, n8587_o, n8572_o, n8562_o, n8555_o, n8527_o, n8501_o, n8497_o, n8493_o, n8450_o, n8447_o, n8435_o, n8432_o, n8426_o, n8422_o, n8395_o, n8393_o, n8388_o, n8386_o, n8368_o, n8349_o, n8343_o, n8325_o, n8323_o, n8316_o, n8314_o, n8305_o, n8286_o, n8268_o, n8264_o, n8215_o, n8212_o, n8166_o, n8164_o, n8144_o, n8127_o, n8124_o, n8075_o, n8072_o, n8021_o, n8018_o, n8015_o};
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8971_o = 1'b1;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8971_o = n8329_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8971_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8971_o = n8307_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8971_o = n7686_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8971_o = n7686_o;
      default: n8971_o = n7686_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n8988_o = 2'b10;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8988_o = 2'b10;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8988_o = 2'b10;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n8816_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8988_o = n8709_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8988_o = 2'b01;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8988_o = 2'b10;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8988_o = 2'b01;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8988_o = 2'b10;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8988_o = 2'b10;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8988_o = 2'b10;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8988_o = 2'b10;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8988_o = 2'b10;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8988_o = 2'b10;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8988_o = 2'b10;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8988_o = 2'b01;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8988_o = 2'b10;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8988_o = n8630_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8988_o = 2'b10;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8988_o = n8584_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8988_o = n7687_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8988_o = n7687_o;
      default: n8988_o = n7687_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n8989_o = n8372_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n8989_o = n8358_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n8989_o = n7688_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n8989_o = n7688_o;
      default: n8989_o = n7688_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9031_o = 2'b10;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9031_o = n7921_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9031_o = n7921_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9031_o = n8934_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9031_o = 2'b01;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9031_o = 2'b01;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9031_o = 2'b01;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9031_o = 2'b01;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9031_o = n7921_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9031_o = n8868_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9031_o = 2'b01;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9031_o = 2'b01;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9031_o = n7921_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9031_o = n8835_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9031_o = n8817_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9031_o = n8803_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9031_o = n8785_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9031_o = n7921_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9031_o = n7921_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9031_o = n7921_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9031_o = n7921_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9031_o = n8711_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9031_o = 2'b01;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9031_o = n8692_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9031_o = 2'b10;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9031_o = 2'b11;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9031_o = 2'b11;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9031_o = 2'b11;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9031_o = 2'b11;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9031_o = 2'b11;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9031_o = 2'b11;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9031_o = 2'b11;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9031_o = 2'b10;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9031_o = 2'b11;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9031_o = 2'b11;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9031_o = 2'b11;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9031_o = 2'b11;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9031_o = n7921_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9031_o = 2'b10;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9031_o = n7921_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9031_o = 2'b11;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9031_o = 2'b10;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9031_o = 2'b10;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9031_o = n7921_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9031_o = 2'b10;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9031_o = 2'b10;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9031_o = n7921_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9031_o = n8542_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9031_o = n8518_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9031_o = n7921_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9031_o = 2'b11;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9031_o = n8461_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9031_o = 2'b01;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9031_o = 2'b01;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9031_o = n7921_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9031_o = 2'b01;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9031_o = n7921_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9031_o = n8403_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9031_o = 2'b01;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9031_o = n7921_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9031_o = 2'b01;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9031_o = n8382_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9031_o = 2'b01;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9031_o = 2'b01;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9031_o = n7921_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9031_o = n7921_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9031_o = 2'b11;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9031_o = n7921_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9031_o = n7921_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9031_o = n8299_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9031_o = n8280_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9031_o = 2'b10;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9031_o = n8252_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9031_o = 2'b11;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9031_o = n8195_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9031_o = 2'b11;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9031_o = n8156_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9031_o = n8138_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9031_o = 2'b10;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9031_o = n8112_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9031_o = n7921_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9031_o = n8054_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9031_o = n7921_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9031_o = 2'b11;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9031_o = n7921_o;
      default: n9031_o = n7921_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9034_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9034_o = n8114_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9034_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9034_o = 1'b0;
      default: n9034_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9037_o = n8338_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9037_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9037_o = 1'b0;
      default: n9037_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9042_o = n8560_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9042_o = n8158_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9042_o = n8115_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9042_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9042_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9042_o = n7690_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9042_o = 1'b1;
      default: n9042_o = n7690_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9044_o = n8198_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9044_o = n8057_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9044_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9044_o = 1'b0;
      default: n9044_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9054_o = 1'b1;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9054_o = n8291_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9054_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9054_o = n8219_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9054_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9054_o = n8201_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9054_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9054_o = n8148_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9054_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9054_o = n8079_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9054_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9054_o = n8060_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9054_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9054_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9054_o = 1'b0;
      default: n9054_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9058_o = n8340_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9058_o = n8320_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9058_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9058_o = n8310_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9058_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9058_o = 1'b0;
      default: n9058_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9076_o = 1'b1;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9076_o = n8713_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9076_o = n8694_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9076_o = 1'b1;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9076_o = 1'b1;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9076_o = 1'b1;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9076_o = 1'b1;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9076_o = 1'b1;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9076_o = 1'b1;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9076_o = 1'b1;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9076_o = 1'b1;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9076_o = 1'b1;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9076_o = 1'b1;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9076_o = 1'b1;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9076_o = 1'b1;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9076_o = 1'b1;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9076_o = 1'b1;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9076_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9076_o = n7701_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9076_o = n7701_o;
      default: n9076_o = n7701_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9078_o = n8640_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9078_o = n8631_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9078_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9078_o = n8000_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9078_o = n8000_o;
      default: n9078_o = n8000_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9081_o = 1'b1;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9081_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9081_o = 1'b0;
      default: n9081_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9084_o = 1'b1;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9084_o = n7894_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9084_o = n7894_o;
      default: n9084_o = n7894_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9087_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9087_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9087_o = 1'b0;
      default: n9087_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9091_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9091_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9091_o = 1'b0;
      default: n9091_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9095_o = n8464_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9095_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9095_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9095_o = 1'b0;
      default: n9095_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9098_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9098_o = n7721_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9098_o = n7721_o;
      default: n9098_o = n7721_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9103_o = 1'b1;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9103_o = 1'b1;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9103_o = 1'b1;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9103_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9103_o = n7923_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9103_o = n7923_o;
      default: n9103_o = n7923_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9105_o = n8466_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9105_o = n8423_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9105_o = n8375_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9105_o = n8361_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9105_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9105_o = 1'b0;
      default: n9105_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9110_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9110_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9110_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9110_o = 1'b0;
      default: n9110_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9113_o = n8469_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9113_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9113_o = 1'b0;
      default: n9113_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9119_o = 1'b1;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9119_o = n8874_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9119_o = n8471_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9119_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9119_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9119_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9119_o = n7727_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9119_o = n7727_o;
      default: n9119_o = n7727_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9123_o = n8937_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9123_o = 1'b1;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9123_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9123_o = n8406_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9123_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9123_o = 1'b0;
      default: n9123_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9128_o = 1'b1;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9128_o = 1'b1;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9128_o = 1'b1;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9128_o = n7963_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9128_o = n7963_o;
      default: n9128_o = n7963_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9129_o = n8961_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9129_o = n8912_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9129_o = n8845_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9129_o = n7734_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9129_o = n7734_o;
      default: n9129_o = n7734_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9133_o = 1'b1;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9133_o = 1'b1;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9133_o = 1'b1;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9133_o = n7738_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9133_o = n7738_o;
      default: n9133_o = n7738_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9136_o = 1'b1;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9136_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9136_o = 1'b0;
      default: n9136_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9140_o = 1'b1;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9140_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9140_o = 1'b0;
      default: n9140_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9142_o = n8766_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9142_o = n7740_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9142_o = n7740_o;
      default: n9142_o = n7740_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9143_o = n8768_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9143_o = n8391_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9143_o = n8003_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9143_o = n8003_o;
      default: n9143_o = n8003_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9146_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9146_o = n8202_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9146_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9146_o = n8061_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9146_o = n2157_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9146_o = n2157_o;
      default: n9146_o = n2157_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9148_o = n8901_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9148_o = 1'b0;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9148_o = 1'b0;
      default: n9148_o = 1'b0;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9150_o = 1'b1;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9150_o = n7785_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9150_o = n7785_o;
      default: n9150_o = n7785_o;
    endcase
  assign n9151_o = n1909_o[20];
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9152_o = 1'b1;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9152_o = 1'b1;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9152_o = n9151_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9152_o = n9151_o;
      default: n9152_o = n9151_o;
    endcase
  assign n9153_o = n1909_o[21];
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9154_o = 1'b1;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9154_o = 1'b1;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9154_o = n9153_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9154_o = n9153_o;
      default: n9154_o = n9153_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9155_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9155_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9155_o = n8062_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9155_o = n2164_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9155_o = n2164_o;
      default: n9155_o = n2164_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9156_o = 1'b1;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9156_o = n7789_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9156_o = n7789_o;
      default: n9156_o = n7789_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9157_o = n8632_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9157_o = n1960_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9157_o = n1960_o;
      default: n9157_o = n1960_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9158_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9158_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9158_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9158_o = n7791_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9158_o = n7791_o;
      default: n9158_o = n7791_o;
    endcase
  assign n9159_o = n1909_o[27];
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9160_o = 1'b1;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9160_o = 1'b1;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9160_o = n8473_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9160_o = n8408_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9160_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9160_o = n9159_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9160_o = n9159_o;
      default: n9160_o = n9159_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9161_o = n8948_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9161_o = n8927_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9161_o = 1'b1;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9161_o = n8875_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9161_o = n8764_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9161_o = 1'b1;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9161_o = 1'b1;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9161_o = n8511_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9161_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9161_o = n8474_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9161_o = n8409_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9161_o = n7795_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9161_o = n7795_o;
      default: n9161_o = n7795_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9162_o = 1'b1;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9162_o = n8679_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9162_o = n7827_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9162_o = n7827_o;
      default: n9162_o = n7827_o;
    endcase
  assign n9163_o = n7797_o[1];
  assign n9164_o = n7779_o[1];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9165_o = n2184_o ? n9163_o : n9164_o;
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9166_o = n8780_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9166_o = n9165_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9166_o = n9165_o;
      default: n9166_o = n9165_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9167_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9167_o = n7967_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9167_o = n7967_o;
      default: n9167_o = n7967_o;
    endcase
  assign n9168_o = n7797_o[3];
  assign n9169_o = n7779_o[3];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9170_o = n2184_o ? n9168_o : n9169_o;
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9171_o = n8821_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9171_o = n8794_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9171_o = 1'b1;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9171_o = n9170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9171_o = n9170_o;
      default: n9171_o = n9170_o;
    endcase
  assign n9172_o = n7797_o[4];
  assign n9173_o = n7779_o[4];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9174_o = n2184_o ? n9172_o : n9173_o;
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9175_o = n8546_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9175_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9175_o = n8478_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9175_o = n8413_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9175_o = n9174_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9175_o = n9174_o;
      default: n9175_o = n9174_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9176_o = n7828_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9176_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9176_o = 1'b1;
      default: n9176_o = n7828_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9177_o = n8714_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9177_o = n8695_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9177_o = 1'b1;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9177_o = 1'b1;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9177_o = 1'b1;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9177_o = n7987_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9177_o = n7987_o;
      default: n9177_o = n7987_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9178_o = 1'b1;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9178_o = 1'b1;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9178_o = 1'b1;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9178_o = 1'b1;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9178_o = 1'b1;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9178_o = 1'b1;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9178_o = 1'b1;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9178_o = 1'b1;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9178_o = 1'b1;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9178_o = 1'b1;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9178_o = 1'b1;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9178_o = 1'b1;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9178_o = 1'b1;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9178_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9178_o = n7971_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9178_o = n7971_o;
      default: n9178_o = n7971_o;
    endcase
  assign n9179_o = n7801_o[3];
  assign n9180_o = n7781_o[3];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9181_o = n2184_o ? n9179_o : n9180_o;
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = n8952_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9182_o = n9181_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9182_o = n9181_o;
      default: n9182_o = n9181_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9183_o = n8602_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9183_o = n8594_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9183_o = n8577_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9183_o = n8567_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9183_o = n7975_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9183_o = n7975_o;
      default: n9183_o = n7975_o;
    endcase
  assign n9184_o = n7801_o[9];
  assign n9185_o = n7781_o[9];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9186_o = n2184_o ? n9184_o : n9185_o;
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9187_o = n8825_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9187_o = n8798_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9187_o = 1'b1;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9187_o = n8550_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9187_o = n8523_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9187_o = n9186_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9187_o = n9186_o;
      default: n9187_o = n9186_o;
    endcase
  assign n9188_o = n7801_o[10];
  assign n9189_o = n7781_o[10];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9190_o = n2184_o ? n9188_o : n9189_o;
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9191_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9191_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9191_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9191_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9191_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9191_o = n9190_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9191_o = n9190_o;
      default: n9191_o = n9190_o;
    endcase
  assign n9192_o = n7801_o[11];
  assign n9193_o = n7781_o[11];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9194_o = n2184_o ? n9192_o : n9193_o;
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9195_o = 1'b1;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9195_o = 1'b1;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9195_o = n9194_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9195_o = n9194_o;
      default: n9195_o = n9194_o;
    endcase
  assign n9196_o = n7801_o[12];
  assign n9197_o = n7781_o[12];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9198_o = n2184_o ? n9196_o : n9197_o;
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9199_o = n8683_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9199_o = 1'b1;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9199_o = n9198_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9199_o = n9198_o;
      default: n9199_o = n9198_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9200_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9200_o = n8479_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9200_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9200_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9200_o = n8159_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9200_o = n8116_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9200_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9200_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9200_o = n2170_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9200_o = 1'b1;
      default: n9200_o = n2170_o;
    endcase
  assign n9201_o = n7803_o[1];
  assign n9202_o = n7601_o[1];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9203_o = n2184_o ? n9201_o : n9202_o;
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9204_o = n8483_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9204_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9204_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9204_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9204_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9204_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9204_o = n8256_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9204_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9204_o = n9203_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9204_o = n9203_o;
      default: n9204_o = n9203_o;
    endcase
  assign n9205_o = n1909_o[67];
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9206_o = n8877_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9206_o = n9205_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9206_o = n9205_o;
      default: n9206_o = n9205_o;
    endcase
  assign n9207_o = n1909_o[68];
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9208_o = n8939_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9208_o = 1'b1;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9208_o = n9207_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9208_o = n9207_o;
      default: n9208_o = n9207_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9209_o = n8551_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9209_o = n7806_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9209_o = n7806_o;
      default: n9209_o = n7806_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9210_o = 1'b1;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9210_o = n8300_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9210_o = n8257_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9210_o = n8203_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9210_o = n8160_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9210_o = n8117_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9210_o = n8063_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9210_o = n7832_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9210_o = n7832_o;
      default: n9210_o = n7832_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9211_o = n8826_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9211_o = 1'b1;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9211_o = n7831_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9211_o = n7831_o;
      default: n9211_o = n7831_o;
    endcase
  assign n9212_o = n7810_o[0];
  assign n9213_o = n7782_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9214_o = n2184_o ? n9212_o : n9213_o;
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9215_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9215_o = n8284_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9215_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9215_o = n8261_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9215_o = n8207_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9215_o = n8142_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9215_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9215_o = n8121_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9215_o = n8067_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9215_o = n9214_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9215_o = n9214_o;
      default: n9215_o = n9214_o;
    endcase
  assign n9216_o = n1909_o[79];
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9217_o = 1'b1;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9217_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9217_o = n9216_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9217_o = n9216_o;
      default: n9217_o = n9216_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9218_o = n8859_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9218_o = n8484_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9218_o = n7815_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9218_o = n7815_o;
      default: n9218_o = n7815_o;
    endcase
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9219_o = n8414_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9219_o = n1925_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9219_o = n1925_o;
      default: n9219_o = n1925_o;
    endcase
  assign n9220_o = n1909_o[84];
  assign n9221_o = n7783_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9222_o = n2184_o ? n9220_o : n9221_o;
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9223_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9223_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9223_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9223_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9223_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9223_o = n9222_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9223_o = n9222_o;
      default: n9223_o = n9222_o;
    endcase
  assign n9224_o = n1909_o[85];
  assign n9225_o = n7783_o[1];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9226_o = n2184_o ? n9224_o : n9225_o;
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9227_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9227_o = n8488_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9227_o = n8418_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9227_o = n9226_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9227_o = n9226_o;
      default: n9227_o = n9226_o;
    endcase
  assign n9228_o = n1909_o[86];
  assign n9229_o = n7783_o[2];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9230_o = n2184_o ? n9228_o : n9229_o;
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9231_o = n8441_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9231_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9231_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9231_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9231_o = n9230_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9231_o = n9230_o;
      default: n9231_o = n9230_o;
    endcase
  assign n9232_o = n1909_o[87];
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9233_o = 1'b1;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9233_o = n9232_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9233_o = n9232_o;
      default: n9233_o = n9232_o;
    endcase
  assign n9234_o = n1909_o[88];
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9235_o = n8379_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9235_o = n8356_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9235_o = n9234_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9235_o = n9234_o;
      default: n9235_o = n9234_o;
    endcase
  assign n9237_o = n1909_o[28];
  assign n9238_o = n7797_o[0];
  assign n9239_o = n7779_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9240_o = n2184_o ? n9238_o : n9239_o;
  assign n9244_o = n7801_o[2];
  assign n9245_o = n7781_o[2];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9246_o = n2184_o ? n9244_o : n9245_o;
  assign n9250_o = n7801_o[8:5];
  assign n9251_o = n7781_o[8:5];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9252_o = n2184_o ? n9250_o : n9251_o;
  assign n9259_o = n7801_o[15:13];
  assign n9260_o = n7781_o[15:13];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9261_o = n2184_o ? n9259_o : n9260_o;
  assign n9262_o = n7803_o[3:2];
  assign n9263_o = n7601_o[3:2];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9264_o = n2184_o ? n9262_o : n9263_o;
  assign n9265_o = n7803_o[0];
  assign n9266_o = n7601_o[0];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9267_o = n2184_o ? n9265_o : n9266_o;
  assign n9269_o = n7810_o[1];
  assign n9270_o = n7782_o[1];
  /* TG68KdotC_Kernel.vhd:1649:17  */
  assign n9271_o = n2184_o ? n9269_o : n9270_o;
  assign n9272_o = n1909_o[78:75];
  assign n9280_o = n7853_o[23];
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n8963_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9281_o = n9280_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9281_o = n9280_o;
      default: n9281_o = n9280_o;
    endcase
  assign n9282_o = n7853_o[25:24];
  assign n9283_o = n7853_o[22:17];
  /* TG68KdotC_Kernel.vhd:3263:25  */
  always @*
    case (n8968_o)
      85'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9329_o = n7937_o;
      85'b0100000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9329_o = n7937_o;
      85'b0010000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9329_o = n7937_o;
      85'b0001000000000000000000000000000000000000000000000000000000000000000000000000000000000: n9329_o = n8941_o;
      85'b0000100000000000000000000000000000000000000000000000000000000000000000000000000000000: n9329_o = n8920_o;
      85'b0000010000000000000000000000000000000000000000000000000000000000000000000000000000000: n9329_o = 7'b1011100;
      85'b0000001000000000000000000000000000000000000000000000000000000000000000000000000000000: n9329_o = n8903_o;
      85'b0000000100000000000000000000000000000000000000000000000000000000000000000000000000000: n9329_o = 7'b1011010;
      85'b0000000010000000000000000000000000000000000000000000000000000000000000000000000000000: n9329_o = n7937_o;
      85'b0000000001000000000000000000000000000000000000000000000000000000000000000000000000000: n9329_o = n8870_o;
      85'b0000000000100000000000000000000000000000000000000000000000000000000000000000000000000: n9329_o = n8853_o;
      85'b0000000000010000000000000000000000000000000000000000000000000000000000000000000000000: n9329_o = 7'b1010110;
      85'b0000000000001000000000000000000000000000000000000000000000000000000000000000000000000: n9329_o = n7937_o;
      85'b0000000000000100000000000000000000000000000000000000000000000000000000000000000000000: n9329_o = 7'b1010010;
      85'b0000000000000010000000000000000000000000000000000000000000000000000000000000000000000: n9329_o = n8828_o;
      85'b0000000000000001000000000000000000000000000000000000000000000000000000000000000000000: n9329_o = 7'b1010000;
      85'b0000000000000000100000000000000000000000000000000000000000000000000000000000000000000: n9329_o = 7'b1001111;
      85'b0000000000000000010000000000000000000000000000000000000000000000000000000000000000000: n9329_o = n7937_o;
      85'b0000000000000000001000000000000000000000000000000000000000000000000000000000000000000: n9329_o = n7937_o;
      85'b0000000000000000000100000000000000000000000000000000000000000000000000000000000000000: n9329_o = 7'b0110001;
      85'b0000000000000000000010000000000000000000000000000000000000000000000000000000000000000: n9329_o = 7'b0000001;
      85'b0000000000000000000001000000000000000000000000000000000000000000000000000000000000000: n9329_o = n8717_o;
      85'b0000000000000000000000100000000000000000000000000000000000000000000000000000000000000: n9329_o = 7'b0101110;
      85'b0000000000000000000000010000000000000000000000000000000000000000000000000000000000000: n9329_o = n8698_o;
      85'b0000000000000000000000001000000000000000000000000000000000000000000000000000000000000: n9329_o = 7'b0101100;
      85'b0000000000000000000000000100000000000000000000000000000000000000000000000000000000000: n9329_o = 7'b0110011;
      85'b0000000000000000000000000010000000000000000000000000000000000000000000000000000000000: n9329_o = 7'b0111101;
      85'b0000000000000000000000000001000000000000000000000000000000000000000000000000000000000: n9329_o = 7'b0111100;
      85'b0000000000000000000000000000100000000000000000000000000000000000000000000000000000000: n9329_o = 7'b0111011;
      85'b0000000000000000000000000000010000000000000000000000000000000000000000000000000000000: n9329_o = 7'b0111010;
      85'b0000000000000000000000000000001000000000000000000000000000000000000000000000000000000: n9329_o = 7'b0111001;
      85'b0000000000000000000000000000000100000000000000000000000000000000000000000000000000000: n9329_o = 7'b0111000;
      85'b0000000000000000000000000000000010000000000000000000000000000000000000000000000000000: n9329_o = 7'b0011000;
      85'b0000000000000000000000000000000001000000000000000000000000000000000000000000000000000: n9329_o = 7'b0110110;
      85'b0000000000000000000000000000000000100000000000000000000000000000000000000000000000000: n9329_o = 7'b0110101;
      85'b0000000000000000000000000000000000010000000000000000000000000000000000000000000000000: n9329_o = n8635_o;
      85'b0000000000000000000000000000000000001000000000000000000000000000000000000000000000000: n9329_o = 7'b0110011;
      85'b0000000000000000000000000000000000000100000000000000000000000000000000000000000000000: n9329_o = n7937_o;
      85'b0000000000000000000000000000000000000010000000000000000000000000000000000000000000000: n9329_o = 7'b0100110;
      85'b0000000000000000000000000000000000000001000000000000000000000000000000000000000000000: n9329_o = n7937_o;
      85'b0000000000000000000000000000000000000000100000000000000000000000000000000000000000000: n9329_o = 7'b0100100;
      85'b0000000000000000000000000000000000000000010000000000000000000000000000000000000000000: n9329_o = n7937_o;
      85'b0000000000000000000000000000000000000000001000000000000000000000000000000000000000000: n9329_o = n7937_o;
      85'b0000000000000000000000000000000000000000000100000000000000000000000000000000000000000: n9329_o = n7937_o;
      85'b0000000000000000000000000000000000000000000010000000000000000000000000000000000000000: n9329_o = 7'b0100000;
      85'b0000000000000000000000000000000000000000000001000000000000000000000000000000000000000: n9329_o = 7'b0011111;
      85'b0000000000000000000000000000000000000000000000100000000000000000000000000000000000000: n9329_o = n7937_o;
      85'b0000000000000000000000000000000000000000000000010000000000000000000000000000000000000: n9329_o = n8553_o;
      85'b0000000000000000000000000000000000000000000000001000000000000000000000000000000000000: n9329_o = n8525_o;
      85'b0000000000000000000000000000000000000000000000000100000000000000000000000000000000000: n9329_o = n7937_o;
      85'b0000000000000000000000000000000000000000000000000010000000000000000000000000000000000: n9329_o = 7'b0011000;
      85'b0000000000000000000000000000000000000000000000000001000000000000000000000000000000000: n9329_o = n8491_o;
      85'b0000000000000000000000000000000000000000000000000000100000000000000000000000000000000: n9329_o = 7'b1000101;
      85'b0000000000000000000000000000000000000000000000000000010000000000000000000000000000000: n9329_o = 7'b1000100;
      85'b0000000000000000000000000000000000000000000000000000001000000000000000000000000000000: n9329_o = 7'b1000011;
      85'b0000000000000000000000000000000000000000000000000000000100000000000000000000000000000: n9329_o = 7'b1000010;
      85'b0000000000000000000000000000000000000000000000000000000010000000000000000000000000000: n9329_o = 7'b1000001;
      85'b0000000000000000000000000000000000000000000000000000000001000000000000000000000000000: n9329_o = n8420_o;
      85'b0000000000000000000000000000000000000000000000000000000000100000000000000000000000000: n9329_o = 7'b0111111;
      85'b0000000000000000000000000000000000000000000000000000000000010000000000000000000000000: n9329_o = n7937_o;
      85'b0000000000000000000000000000000000000000000000000000000000001000000000000000000000000: n9329_o = 7'b1001100;
      85'b0000000000000000000000000000000000000000000000000000000000000100000000000000000000000: n9329_o = n8384_o;
      85'b0000000000000000000000000000000000000000000000000000000000000010000000000000000000000: n9329_o = 7'b1001010;
      85'b0000000000000000000000000000000000000000000000000000000000000001000000000000000000000: n9329_o = 7'b1001001;
      85'b0000000000000000000000000000000000000000000000000000000000000000100000000000000000000: n9329_o = n8334_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000010000000000000000000: n9329_o = 7'b0000001;
      85'b0000000000000000000000000000000000000000000000000000000000000000001000000000000000000: n9329_o = 7'b0011000;
      85'b0000000000000000000000000000000000000000000000000000000000000000000100000000000000000: n9329_o = 7'b0000001;
      85'b0000000000000000000000000000000000000000000000000000000000000000000010000000000000000: n9329_o = n8312_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000001000000000000000: n9329_o = n8303_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000100000000000000: n9329_o = 7'b0010010;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000010000000000000: n9329_o = 7'b0010001;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000001000000000000: n9329_o = n8262_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000100000000000: n9329_o = 7'b0000001;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000010000000000: n9329_o = n8210_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000001000000000: n9329_o = 7'b0000001;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000100000000: n9329_o = n8162_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000010000000: n9329_o = 7'b0001110;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000001000000: n9329_o = 7'b0001101;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000100000: n9329_o = n8122_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000010000: n9329_o = n7937_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000001000: n9329_o = n8070_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000100: n9329_o = n7937_o;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000010: n9329_o = 7'b0000001;
      85'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000001: n9329_o = n7937_o;
      default: n9329_o = n7937_o;
    endcase
  /* TG68KdotC_Kernel.vhd:4049:41  */
  assign n9334_o = exec[33];
  /* TG68KdotC_Kernel.vhd:4049:33  */
  assign n9335_o = n9334_o & clkena_lw;
  /* TG68KdotC_Kernel.vhd:4050:27  */
  assign n9336_o = brief[11:0];
  /* TG68KdotC_Kernel.vhd:4051:47  */
  assign n9337_o = reg_qa[2:0];
  /* TG68KdotC_Kernel.vhd:4051:19  */
  assign n9339_o = n9336_o == 12'b000000000000;
  /* TG68KdotC_Kernel.vhd:4052:47  */
  assign n9340_o = reg_qa[2:0];
  /* TG68KdotC_Kernel.vhd:4052:19  */
  assign n9342_o = n9336_o == 12'b000000000001;
  /* TG68KdotC_Kernel.vhd:4053:48  */
  assign n9343_o = reg_qa[3:0];
  /* TG68KdotC_Kernel.vhd:4053:19  */
  assign n9345_o = n9336_o == 12'b000000000010;
  /* TG68KdotC_Kernel.vhd:4054:19  */
  assign n9347_o = n9336_o == 12'b100000000000;
  /* TG68KdotC_Kernel.vhd:4055:19  */
  assign n9349_o = n9336_o == 12'b100000000001;
  /* TG68KdotC_Kernel.vhd:4056:19  */
  assign n9351_o = n9336_o == 12'b100000000010;
  /* TG68KdotC_Kernel.vhd:4057:19  */
  assign n9353_o = n9336_o == 12'b100000000011;
  /* TG68KdotC_Kernel.vhd:4058:19  */
  assign n9355_o = n9336_o == 12'b100000000100;
  assign n9356_o = {n9355_o, n9353_o, n9351_o, n9349_o, n9347_o, n9345_o, n9342_o, n9339_o};
  /* TG68KdotC_Kernel.vhd:4050:17  */
  always @*
    case (n9356_o)
      8'b10000000: n9357_o = vbr;
      8'b01000000: n9357_o = vbr;
      8'b00100000: n9357_o = vbr;
      8'b00010000: n9357_o = reg_qa;
      8'b00001000: n9357_o = vbr;
      8'b00000100: n9357_o = vbr;
      8'b00000010: n9357_o = vbr;
      8'b00000001: n9357_o = vbr;
      default: n9357_o = vbr;
    endcase
  /* TG68KdotC_Kernel.vhd:4050:17  */
  always @*
    case (n9356_o)
      8'b10000000: n9358_o = cacr;
      8'b01000000: n9358_o = cacr;
      8'b00100000: n9358_o = cacr;
      8'b00010000: n9358_o = cacr;
      8'b00001000: n9358_o = cacr;
      8'b00000100: n9358_o = n9343_o;
      8'b00000010: n9358_o = cacr;
      8'b00000001: n9358_o = cacr;
      default: n9358_o = cacr;
    endcase
  /* TG68KdotC_Kernel.vhd:4050:17  */
  always @*
    case (n9356_o)
      8'b10000000: n9359_o = dfc;
      8'b01000000: n9359_o = dfc;
      8'b00100000: n9359_o = dfc;
      8'b00010000: n9359_o = dfc;
      8'b00001000: n9359_o = dfc;
      8'b00000100: n9359_o = dfc;
      8'b00000010: n9359_o = n9340_o;
      8'b00000001: n9359_o = dfc;
      default: n9359_o = dfc;
    endcase
  /* TG68KdotC_Kernel.vhd:4050:17  */
  always @*
    case (n9356_o)
      8'b10000000: n9360_o = sfc;
      8'b01000000: n9360_o = sfc;
      8'b00100000: n9360_o = sfc;
      8'b00010000: n9360_o = sfc;
      8'b00001000: n9360_o = sfc;
      8'b00000100: n9360_o = sfc;
      8'b00000010: n9360_o = sfc;
      8'b00000001: n9360_o = n9337_o;
      default: n9360_o = sfc;
    endcase
  /* TG68KdotC_Kernel.vhd:4049:11  */
  assign n9361_o = n9335_o ? n9357_o : vbr;
  /* TG68KdotC_Kernel.vhd:4049:11  */
  assign n9362_o = n9335_o ? n9358_o : cacr;
  /* TG68KdotC_Kernel.vhd:4049:11  */
  assign n9363_o = n9335_o ? n9359_o : dfc;
  /* TG68KdotC_Kernel.vhd:4049:11  */
  assign n9364_o = n9335_o ? n9360_o : sfc;
  /* TG68KdotC_Kernel.vhd:4046:11  */
  assign n9366_o = reset ? 32'b00000000000000000000000000000000 : n9361_o;
  /* TG68KdotC_Kernel.vhd:4046:11  */
  assign n9368_o = reset ? 4'b0000 : n9362_o;
  /* TG68KdotC_Kernel.vhd:4046:11  */
  assign n9369_o = reset ? dfc : n9363_o;
  /* TG68KdotC_Kernel.vhd:4046:11  */
  assign n9370_o = reset ? sfc : n9364_o;
  /* TG68KdotC_Kernel.vhd:4065:19  */
  assign n9375_o = brief[11:0];
  /* TG68KdotC_Kernel.vhd:4066:78  */
  assign n9377_o = {29'b00000000000000000000000000000, sfc};
  /* TG68KdotC_Kernel.vhd:4066:17  */
  assign n9379_o = n9375_o == 12'b000000000000;
  /* TG68KdotC_Kernel.vhd:4067:78  */
  assign n9381_o = {29'b00000000000000000000000000000, dfc};
  /* TG68KdotC_Kernel.vhd:4067:17  */
  assign n9383_o = n9375_o == 12'b000000000001;
  /* TG68KdotC_Kernel.vhd:4068:79  */
  assign n9385_o = cacr & 4'b0011;
  /* TG68KdotC_Kernel.vhd:4068:71  */
  assign n9387_o = {28'b0000000000000000000000000000, n9385_o};
  /* TG68KdotC_Kernel.vhd:4068:11  */
  assign n9389_o = n9375_o == 12'b000000000010;
  /* TG68KdotC_Kernel.vhd:4070:11  */
  assign n9391_o = n9375_o == 12'b100000000001;
  assign n9392_o = {n9391_o, n9389_o, n9383_o, n9379_o};
  /* TG68KdotC_Kernel.vhd:4065:9  */
  always @*
    case (n9392_o)
      4'b1000: n9394_o = vbr;
      4'b0100: n9394_o = n9387_o;
      4'b0010: n9394_o = n9381_o;
      4'b0001: n9394_o = n9377_o;
      default: n9394_o = 32'b00000000000000000000000000000000;
    endcase
  /* TG68KdotC_Kernel.vhd:4084:32  */
  assign n9399_o = exe_opcode[11:8];
  /* TG68KdotC_Kernel.vhd:4085:25  */
  assign n9401_o = n9399_o == 4'b0000;
  /* TG68KdotC_Kernel.vhd:4086:25  */
  assign n9403_o = n9399_o == 4'b0001;
  /* TG68KdotC_Kernel.vhd:4087:65  */
  assign n9404_o = flags[0];
  /* TG68KdotC_Kernel.vhd:4087:56  */
  assign n9405_o = ~n9404_o;
  /* TG68KdotC_Kernel.vhd:4087:82  */
  assign n9406_o = flags[2];
  /* TG68KdotC_Kernel.vhd:4087:73  */
  assign n9407_o = ~n9406_o;
  /* TG68KdotC_Kernel.vhd:4087:69  */
  assign n9408_o = n9405_o & n9407_o;
  /* TG68KdotC_Kernel.vhd:4087:25  */
  assign n9410_o = n9399_o == 4'b0010;
  /* TG68KdotC_Kernel.vhd:4088:60  */
  assign n9411_o = flags[0];
  /* TG68KdotC_Kernel.vhd:4088:72  */
  assign n9412_o = flags[2];
  /* TG68KdotC_Kernel.vhd:4088:64  */
  assign n9413_o = n9411_o | n9412_o;
  /* TG68KdotC_Kernel.vhd:4088:25  */
  assign n9415_o = n9399_o == 4'b0011;
  /* TG68KdotC_Kernel.vhd:4089:64  */
  assign n9416_o = flags[0];
  /* TG68KdotC_Kernel.vhd:4089:55  */
  assign n9417_o = ~n9416_o;
  /* TG68KdotC_Kernel.vhd:4089:25  */
  assign n9419_o = n9399_o == 4'b0100;
  /* TG68KdotC_Kernel.vhd:4090:60  */
  assign n9420_o = flags[0];
  /* TG68KdotC_Kernel.vhd:4090:25  */
  assign n9422_o = n9399_o == 4'b0101;
  /* TG68KdotC_Kernel.vhd:4091:64  */
  assign n9423_o = flags[2];
  /* TG68KdotC_Kernel.vhd:4091:55  */
  assign n9424_o = ~n9423_o;
  /* TG68KdotC_Kernel.vhd:4091:25  */
  assign n9426_o = n9399_o == 4'b0110;
  /* TG68KdotC_Kernel.vhd:4092:60  */
  assign n9427_o = flags[2];
  /* TG68KdotC_Kernel.vhd:4092:25  */
  assign n9429_o = n9399_o == 4'b0111;
  /* TG68KdotC_Kernel.vhd:4093:64  */
  assign n9430_o = flags[1];
  /* TG68KdotC_Kernel.vhd:4093:55  */
  assign n9431_o = ~n9430_o;
  /* TG68KdotC_Kernel.vhd:4093:25  */
  assign n9433_o = n9399_o == 4'b1000;
  /* TG68KdotC_Kernel.vhd:4094:60  */
  assign n9434_o = flags[1];
  /* TG68KdotC_Kernel.vhd:4094:25  */
  assign n9436_o = n9399_o == 4'b1001;
  /* TG68KdotC_Kernel.vhd:4095:64  */
  assign n9437_o = flags[3];
  /* TG68KdotC_Kernel.vhd:4095:55  */
  assign n9438_o = ~n9437_o;
  /* TG68KdotC_Kernel.vhd:4095:25  */
  assign n9440_o = n9399_o == 4'b1010;
  /* TG68KdotC_Kernel.vhd:4096:60  */
  assign n9441_o = flags[3];
  /* TG68KdotC_Kernel.vhd:4096:25  */
  assign n9443_o = n9399_o == 4'b1011;
  /* TG68KdotC_Kernel.vhd:4097:61  */
  assign n9444_o = flags[3];
  /* TG68KdotC_Kernel.vhd:4097:74  */
  assign n9445_o = flags[1];
  /* TG68KdotC_Kernel.vhd:4097:65  */
  assign n9446_o = n9444_o & n9445_o;
  /* TG68KdotC_Kernel.vhd:4097:92  */
  assign n9447_o = flags[3];
  /* TG68KdotC_Kernel.vhd:4097:83  */
  assign n9448_o = ~n9447_o;
  /* TG68KdotC_Kernel.vhd:4097:109  */
  assign n9449_o = flags[1];
  /* TG68KdotC_Kernel.vhd:4097:100  */
  assign n9450_o = ~n9449_o;
  /* TG68KdotC_Kernel.vhd:4097:96  */
  assign n9451_o = n9448_o & n9450_o;
  /* TG68KdotC_Kernel.vhd:4097:79  */
  assign n9452_o = n9446_o | n9451_o;
  /* TG68KdotC_Kernel.vhd:4097:25  */
  assign n9454_o = n9399_o == 4'b1100;
  /* TG68KdotC_Kernel.vhd:4098:61  */
  assign n9455_o = flags[3];
  /* TG68KdotC_Kernel.vhd:4098:78  */
  assign n9456_o = flags[1];
  /* TG68KdotC_Kernel.vhd:4098:69  */
  assign n9457_o = ~n9456_o;
  /* TG68KdotC_Kernel.vhd:4098:65  */
  assign n9458_o = n9455_o & n9457_o;
  /* TG68KdotC_Kernel.vhd:4098:96  */
  assign n9459_o = flags[3];
  /* TG68KdotC_Kernel.vhd:4098:87  */
  assign n9460_o = ~n9459_o;
  /* TG68KdotC_Kernel.vhd:4098:109  */
  assign n9461_o = flags[1];
  /* TG68KdotC_Kernel.vhd:4098:100  */
  assign n9462_o = n9460_o & n9461_o;
  /* TG68KdotC_Kernel.vhd:4098:83  */
  assign n9463_o = n9458_o | n9462_o;
  /* TG68KdotC_Kernel.vhd:4098:25  */
  assign n9465_o = n9399_o == 4'b1101;
  /* TG68KdotC_Kernel.vhd:4099:61  */
  assign n9466_o = flags[3];
  /* TG68KdotC_Kernel.vhd:4099:74  */
  assign n9467_o = flags[1];
  /* TG68KdotC_Kernel.vhd:4099:65  */
  assign n9468_o = n9466_o & n9467_o;
  /* TG68KdotC_Kernel.vhd:4099:91  */
  assign n9469_o = flags[2];
  /* TG68KdotC_Kernel.vhd:4099:82  */
  assign n9470_o = ~n9469_o;
  /* TG68KdotC_Kernel.vhd:4099:78  */
  assign n9471_o = n9468_o & n9470_o;
  /* TG68KdotC_Kernel.vhd:4099:109  */
  assign n9472_o = flags[3];
  /* TG68KdotC_Kernel.vhd:4099:100  */
  assign n9473_o = ~n9472_o;
  /* TG68KdotC_Kernel.vhd:4099:126  */
  assign n9474_o = flags[1];
  /* TG68KdotC_Kernel.vhd:4099:117  */
  assign n9475_o = ~n9474_o;
  /* TG68KdotC_Kernel.vhd:4099:113  */
  assign n9476_o = n9473_o & n9475_o;
  /* TG68KdotC_Kernel.vhd:4099:143  */
  assign n9477_o = flags[2];
  /* TG68KdotC_Kernel.vhd:4099:134  */
  assign n9478_o = ~n9477_o;
  /* TG68KdotC_Kernel.vhd:4099:130  */
  assign n9479_o = n9476_o & n9478_o;
  /* TG68KdotC_Kernel.vhd:4099:96  */
  assign n9480_o = n9471_o | n9479_o;
  /* TG68KdotC_Kernel.vhd:4099:25  */
  assign n9482_o = n9399_o == 4'b1110;
  /* TG68KdotC_Kernel.vhd:4100:61  */
  assign n9483_o = flags[3];
  /* TG68KdotC_Kernel.vhd:4100:78  */
  assign n9484_o = flags[1];
  /* TG68KdotC_Kernel.vhd:4100:69  */
  assign n9485_o = ~n9484_o;
  /* TG68KdotC_Kernel.vhd:4100:65  */
  assign n9486_o = n9483_o & n9485_o;
  /* TG68KdotC_Kernel.vhd:4100:96  */
  assign n9487_o = flags[3];
  /* TG68KdotC_Kernel.vhd:4100:87  */
  assign n9488_o = ~n9487_o;
  /* TG68KdotC_Kernel.vhd:4100:109  */
  assign n9489_o = flags[1];
  /* TG68KdotC_Kernel.vhd:4100:100  */
  assign n9490_o = n9488_o & n9489_o;
  /* TG68KdotC_Kernel.vhd:4100:83  */
  assign n9491_o = n9486_o | n9490_o;
  /* TG68KdotC_Kernel.vhd:4100:122  */
  assign n9492_o = flags[2];
  /* TG68KdotC_Kernel.vhd:4100:114  */
  assign n9493_o = n9491_o | n9492_o;
  /* TG68KdotC_Kernel.vhd:4100:25  */
  assign n9495_o = n9399_o == 4'b1111;
  assign n9496_o = {n9495_o, n9482_o, n9465_o, n9454_o, n9443_o, n9440_o, n9436_o, n9433_o, n9429_o, n9426_o, n9422_o, n9419_o, n9415_o, n9410_o, n9403_o, n9401_o};
  /* TG68KdotC_Kernel.vhd:4084:17  */
  always @*
    case (n9496_o)
      16'b1000000000000000: n9499_o = n9493_o;
      16'b0100000000000000: n9499_o = n9480_o;
      16'b0010000000000000: n9499_o = n9463_o;
      16'b0001000000000000: n9499_o = n9452_o;
      16'b0000100000000000: n9499_o = n9441_o;
      16'b0000010000000000: n9499_o = n9438_o;
      16'b0000001000000000: n9499_o = n9434_o;
      16'b0000000100000000: n9499_o = n9431_o;
      16'b0000000010000000: n9499_o = n9427_o;
      16'b0000000001000000: n9499_o = n9424_o;
      16'b0000000000100000: n9499_o = n9420_o;
      16'b0000000000010000: n9499_o = n9417_o;
      16'b0000000000001000: n9499_o = n9413_o;
      16'b0000000000000100: n9499_o = n9408_o;
      16'b0000000000000010: n9499_o = 1'b0;
      16'b0000000000000001: n9499_o = 1'b1;
      default: n9499_o = exe_condition;
    endcase
  /* TG68KdotC_Kernel.vhd:4112:54  */
  assign n9504_o = exec[69];
  /* TG68KdotC_Kernel.vhd:4114:60  */
  assign n9505_o = data_read[15:0];
  /* TG68KdotC_Kernel.vhd:4115:43  */
  assign n9506_o = exec[69];
  /* TG68KdotC_Kernel.vhd:4115:68  */
  assign n9507_o = set[69];
  /* TG68KdotC_Kernel.vhd:4115:62  */
  assign n9508_o = n9506_o | n9507_o;
  /* TG68KdotC_Kernel.vhd:4117:49  */
  assign n9511_o = movem_regaddr == 4'b0000;
  /* TG68KdotC_Kernel.vhd:4118:49  */
  assign n9514_o = movem_regaddr == 4'b0001;
  /* TG68KdotC_Kernel.vhd:4119:49  */
  assign n9517_o = movem_regaddr == 4'b0010;
  /* TG68KdotC_Kernel.vhd:4120:49  */
  assign n9520_o = movem_regaddr == 4'b0011;
  /* TG68KdotC_Kernel.vhd:4121:49  */
  assign n9523_o = movem_regaddr == 4'b0100;
  /* TG68KdotC_Kernel.vhd:4122:49  */
  assign n9526_o = movem_regaddr == 4'b0101;
  /* TG68KdotC_Kernel.vhd:4123:49  */
  assign n9529_o = movem_regaddr == 4'b0110;
  /* TG68KdotC_Kernel.vhd:4124:49  */
  assign n9532_o = movem_regaddr == 4'b0111;
  /* TG68KdotC_Kernel.vhd:4125:49  */
  assign n9535_o = movem_regaddr == 4'b1000;
  /* TG68KdotC_Kernel.vhd:4126:49  */
  assign n9538_o = movem_regaddr == 4'b1001;
  /* TG68KdotC_Kernel.vhd:4127:49  */
  assign n9541_o = movem_regaddr == 4'b1010;
  /* TG68KdotC_Kernel.vhd:4128:49  */
  assign n9544_o = movem_regaddr == 4'b1011;
  /* TG68KdotC_Kernel.vhd:4129:49  */
  assign n9547_o = movem_regaddr == 4'b1100;
  /* TG68KdotC_Kernel.vhd:4130:49  */
  assign n9550_o = movem_regaddr == 4'b1101;
  /* TG68KdotC_Kernel.vhd:4131:49  */
  assign n9553_o = movem_regaddr == 4'b1110;
  /* TG68KdotC_Kernel.vhd:4132:49  */
  assign n9556_o = movem_regaddr == 4'b1111;
  assign n9557_o = {n9556_o, n9553_o, n9550_o, n9547_o, n9544_o, n9541_o, n9538_o, n9535_o, n9532_o, n9529_o, n9526_o, n9523_o, n9520_o, n9517_o, n9514_o, n9511_o};
  assign n9558_o = sndopc[0];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9557_o)
      16'b1000000000000000: n9559_o = n9558_o;
      16'b0100000000000000: n9559_o = n9558_o;
      16'b0010000000000000: n9559_o = n9558_o;
      16'b0001000000000000: n9559_o = n9558_o;
      16'b0000100000000000: n9559_o = n9558_o;
      16'b0000010000000000: n9559_o = n9558_o;
      16'b0000001000000000: n9559_o = n9558_o;
      16'b0000000100000000: n9559_o = n9558_o;
      16'b0000000010000000: n9559_o = n9558_o;
      16'b0000000001000000: n9559_o = n9558_o;
      16'b0000000000100000: n9559_o = n9558_o;
      16'b0000000000010000: n9559_o = n9558_o;
      16'b0000000000001000: n9559_o = n9558_o;
      16'b0000000000000100: n9559_o = n9558_o;
      16'b0000000000000010: n9559_o = n9558_o;
      16'b0000000000000001: n9559_o = 1'b0;
      default: n9559_o = n9558_o;
    endcase
  assign n9560_o = sndopc[1];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9557_o)
      16'b1000000000000000: n9561_o = n9560_o;
      16'b0100000000000000: n9561_o = n9560_o;
      16'b0010000000000000: n9561_o = n9560_o;
      16'b0001000000000000: n9561_o = n9560_o;
      16'b0000100000000000: n9561_o = n9560_o;
      16'b0000010000000000: n9561_o = n9560_o;
      16'b0000001000000000: n9561_o = n9560_o;
      16'b0000000100000000: n9561_o = n9560_o;
      16'b0000000010000000: n9561_o = n9560_o;
      16'b0000000001000000: n9561_o = n9560_o;
      16'b0000000000100000: n9561_o = n9560_o;
      16'b0000000000010000: n9561_o = n9560_o;
      16'b0000000000001000: n9561_o = n9560_o;
      16'b0000000000000100: n9561_o = n9560_o;
      16'b0000000000000010: n9561_o = 1'b0;
      16'b0000000000000001: n9561_o = n9560_o;
      default: n9561_o = n9560_o;
    endcase
  assign n9562_o = sndopc[2];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9557_o)
      16'b1000000000000000: n9563_o = n9562_o;
      16'b0100000000000000: n9563_o = n9562_o;
      16'b0010000000000000: n9563_o = n9562_o;
      16'b0001000000000000: n9563_o = n9562_o;
      16'b0000100000000000: n9563_o = n9562_o;
      16'b0000010000000000: n9563_o = n9562_o;
      16'b0000001000000000: n9563_o = n9562_o;
      16'b0000000100000000: n9563_o = n9562_o;
      16'b0000000010000000: n9563_o = n9562_o;
      16'b0000000001000000: n9563_o = n9562_o;
      16'b0000000000100000: n9563_o = n9562_o;
      16'b0000000000010000: n9563_o = n9562_o;
      16'b0000000000001000: n9563_o = n9562_o;
      16'b0000000000000100: n9563_o = 1'b0;
      16'b0000000000000010: n9563_o = n9562_o;
      16'b0000000000000001: n9563_o = n9562_o;
      default: n9563_o = n9562_o;
    endcase
  assign n9564_o = sndopc[3];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9557_o)
      16'b1000000000000000: n9565_o = n9564_o;
      16'b0100000000000000: n9565_o = n9564_o;
      16'b0010000000000000: n9565_o = n9564_o;
      16'b0001000000000000: n9565_o = n9564_o;
      16'b0000100000000000: n9565_o = n9564_o;
      16'b0000010000000000: n9565_o = n9564_o;
      16'b0000001000000000: n9565_o = n9564_o;
      16'b0000000100000000: n9565_o = n9564_o;
      16'b0000000010000000: n9565_o = n9564_o;
      16'b0000000001000000: n9565_o = n9564_o;
      16'b0000000000100000: n9565_o = n9564_o;
      16'b0000000000010000: n9565_o = n9564_o;
      16'b0000000000001000: n9565_o = 1'b0;
      16'b0000000000000100: n9565_o = n9564_o;
      16'b0000000000000010: n9565_o = n9564_o;
      16'b0000000000000001: n9565_o = n9564_o;
      default: n9565_o = n9564_o;
    endcase
  assign n9566_o = sndopc[4];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9557_o)
      16'b1000000000000000: n9567_o = n9566_o;
      16'b0100000000000000: n9567_o = n9566_o;
      16'b0010000000000000: n9567_o = n9566_o;
      16'b0001000000000000: n9567_o = n9566_o;
      16'b0000100000000000: n9567_o = n9566_o;
      16'b0000010000000000: n9567_o = n9566_o;
      16'b0000001000000000: n9567_o = n9566_o;
      16'b0000000100000000: n9567_o = n9566_o;
      16'b0000000010000000: n9567_o = n9566_o;
      16'b0000000001000000: n9567_o = n9566_o;
      16'b0000000000100000: n9567_o = n9566_o;
      16'b0000000000010000: n9567_o = 1'b0;
      16'b0000000000001000: n9567_o = n9566_o;
      16'b0000000000000100: n9567_o = n9566_o;
      16'b0000000000000010: n9567_o = n9566_o;
      16'b0000000000000001: n9567_o = n9566_o;
      default: n9567_o = n9566_o;
    endcase
  assign n9568_o = sndopc[5];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9557_o)
      16'b1000000000000000: n9569_o = n9568_o;
      16'b0100000000000000: n9569_o = n9568_o;
      16'b0010000000000000: n9569_o = n9568_o;
      16'b0001000000000000: n9569_o = n9568_o;
      16'b0000100000000000: n9569_o = n9568_o;
      16'b0000010000000000: n9569_o = n9568_o;
      16'b0000001000000000: n9569_o = n9568_o;
      16'b0000000100000000: n9569_o = n9568_o;
      16'b0000000010000000: n9569_o = n9568_o;
      16'b0000000001000000: n9569_o = n9568_o;
      16'b0000000000100000: n9569_o = 1'b0;
      16'b0000000000010000: n9569_o = n9568_o;
      16'b0000000000001000: n9569_o = n9568_o;
      16'b0000000000000100: n9569_o = n9568_o;
      16'b0000000000000010: n9569_o = n9568_o;
      16'b0000000000000001: n9569_o = n9568_o;
      default: n9569_o = n9568_o;
    endcase
  assign n9570_o = sndopc[6];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9557_o)
      16'b1000000000000000: n9571_o = n9570_o;
      16'b0100000000000000: n9571_o = n9570_o;
      16'b0010000000000000: n9571_o = n9570_o;
      16'b0001000000000000: n9571_o = n9570_o;
      16'b0000100000000000: n9571_o = n9570_o;
      16'b0000010000000000: n9571_o = n9570_o;
      16'b0000001000000000: n9571_o = n9570_o;
      16'b0000000100000000: n9571_o = n9570_o;
      16'b0000000010000000: n9571_o = n9570_o;
      16'b0000000001000000: n9571_o = 1'b0;
      16'b0000000000100000: n9571_o = n9570_o;
      16'b0000000000010000: n9571_o = n9570_o;
      16'b0000000000001000: n9571_o = n9570_o;
      16'b0000000000000100: n9571_o = n9570_o;
      16'b0000000000000010: n9571_o = n9570_o;
      16'b0000000000000001: n9571_o = n9570_o;
      default: n9571_o = n9570_o;
    endcase
  assign n9572_o = sndopc[7];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9557_o)
      16'b1000000000000000: n9573_o = n9572_o;
      16'b0100000000000000: n9573_o = n9572_o;
      16'b0010000000000000: n9573_o = n9572_o;
      16'b0001000000000000: n9573_o = n9572_o;
      16'b0000100000000000: n9573_o = n9572_o;
      16'b0000010000000000: n9573_o = n9572_o;
      16'b0000001000000000: n9573_o = n9572_o;
      16'b0000000100000000: n9573_o = n9572_o;
      16'b0000000010000000: n9573_o = 1'b0;
      16'b0000000001000000: n9573_o = n9572_o;
      16'b0000000000100000: n9573_o = n9572_o;
      16'b0000000000010000: n9573_o = n9572_o;
      16'b0000000000001000: n9573_o = n9572_o;
      16'b0000000000000100: n9573_o = n9572_o;
      16'b0000000000000010: n9573_o = n9572_o;
      16'b0000000000000001: n9573_o = n9572_o;
      default: n9573_o = n9572_o;
    endcase
  assign n9574_o = sndopc[8];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9557_o)
      16'b1000000000000000: n9575_o = n9574_o;
      16'b0100000000000000: n9575_o = n9574_o;
      16'b0010000000000000: n9575_o = n9574_o;
      16'b0001000000000000: n9575_o = n9574_o;
      16'b0000100000000000: n9575_o = n9574_o;
      16'b0000010000000000: n9575_o = n9574_o;
      16'b0000001000000000: n9575_o = n9574_o;
      16'b0000000100000000: n9575_o = 1'b0;
      16'b0000000010000000: n9575_o = n9574_o;
      16'b0000000001000000: n9575_o = n9574_o;
      16'b0000000000100000: n9575_o = n9574_o;
      16'b0000000000010000: n9575_o = n9574_o;
      16'b0000000000001000: n9575_o = n9574_o;
      16'b0000000000000100: n9575_o = n9574_o;
      16'b0000000000000010: n9575_o = n9574_o;
      16'b0000000000000001: n9575_o = n9574_o;
      default: n9575_o = n9574_o;
    endcase
  assign n9576_o = sndopc[9];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9557_o)
      16'b1000000000000000: n9577_o = n9576_o;
      16'b0100000000000000: n9577_o = n9576_o;
      16'b0010000000000000: n9577_o = n9576_o;
      16'b0001000000000000: n9577_o = n9576_o;
      16'b0000100000000000: n9577_o = n9576_o;
      16'b0000010000000000: n9577_o = n9576_o;
      16'b0000001000000000: n9577_o = 1'b0;
      16'b0000000100000000: n9577_o = n9576_o;
      16'b0000000010000000: n9577_o = n9576_o;
      16'b0000000001000000: n9577_o = n9576_o;
      16'b0000000000100000: n9577_o = n9576_o;
      16'b0000000000010000: n9577_o = n9576_o;
      16'b0000000000001000: n9577_o = n9576_o;
      16'b0000000000000100: n9577_o = n9576_o;
      16'b0000000000000010: n9577_o = n9576_o;
      16'b0000000000000001: n9577_o = n9576_o;
      default: n9577_o = n9576_o;
    endcase
  assign n9578_o = sndopc[10];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9557_o)
      16'b1000000000000000: n9579_o = n9578_o;
      16'b0100000000000000: n9579_o = n9578_o;
      16'b0010000000000000: n9579_o = n9578_o;
      16'b0001000000000000: n9579_o = n9578_o;
      16'b0000100000000000: n9579_o = n9578_o;
      16'b0000010000000000: n9579_o = 1'b0;
      16'b0000001000000000: n9579_o = n9578_o;
      16'b0000000100000000: n9579_o = n9578_o;
      16'b0000000010000000: n9579_o = n9578_o;
      16'b0000000001000000: n9579_o = n9578_o;
      16'b0000000000100000: n9579_o = n9578_o;
      16'b0000000000010000: n9579_o = n9578_o;
      16'b0000000000001000: n9579_o = n9578_o;
      16'b0000000000000100: n9579_o = n9578_o;
      16'b0000000000000010: n9579_o = n9578_o;
      16'b0000000000000001: n9579_o = n9578_o;
      default: n9579_o = n9578_o;
    endcase
  assign n9580_o = sndopc[11];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9557_o)
      16'b1000000000000000: n9581_o = n9580_o;
      16'b0100000000000000: n9581_o = n9580_o;
      16'b0010000000000000: n9581_o = n9580_o;
      16'b0001000000000000: n9581_o = n9580_o;
      16'b0000100000000000: n9581_o = 1'b0;
      16'b0000010000000000: n9581_o = n9580_o;
      16'b0000001000000000: n9581_o = n9580_o;
      16'b0000000100000000: n9581_o = n9580_o;
      16'b0000000010000000: n9581_o = n9580_o;
      16'b0000000001000000: n9581_o = n9580_o;
      16'b0000000000100000: n9581_o = n9580_o;
      16'b0000000000010000: n9581_o = n9580_o;
      16'b0000000000001000: n9581_o = n9580_o;
      16'b0000000000000100: n9581_o = n9580_o;
      16'b0000000000000010: n9581_o = n9580_o;
      16'b0000000000000001: n9581_o = n9580_o;
      default: n9581_o = n9580_o;
    endcase
  assign n9582_o = sndopc[12];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9557_o)
      16'b1000000000000000: n9583_o = n9582_o;
      16'b0100000000000000: n9583_o = n9582_o;
      16'b0010000000000000: n9583_o = n9582_o;
      16'b0001000000000000: n9583_o = 1'b0;
      16'b0000100000000000: n9583_o = n9582_o;
      16'b0000010000000000: n9583_o = n9582_o;
      16'b0000001000000000: n9583_o = n9582_o;
      16'b0000000100000000: n9583_o = n9582_o;
      16'b0000000010000000: n9583_o = n9582_o;
      16'b0000000001000000: n9583_o = n9582_o;
      16'b0000000000100000: n9583_o = n9582_o;
      16'b0000000000010000: n9583_o = n9582_o;
      16'b0000000000001000: n9583_o = n9582_o;
      16'b0000000000000100: n9583_o = n9582_o;
      16'b0000000000000010: n9583_o = n9582_o;
      16'b0000000000000001: n9583_o = n9582_o;
      default: n9583_o = n9582_o;
    endcase
  assign n9584_o = sndopc[13];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9557_o)
      16'b1000000000000000: n9585_o = n9584_o;
      16'b0100000000000000: n9585_o = n9584_o;
      16'b0010000000000000: n9585_o = 1'b0;
      16'b0001000000000000: n9585_o = n9584_o;
      16'b0000100000000000: n9585_o = n9584_o;
      16'b0000010000000000: n9585_o = n9584_o;
      16'b0000001000000000: n9585_o = n9584_o;
      16'b0000000100000000: n9585_o = n9584_o;
      16'b0000000010000000: n9585_o = n9584_o;
      16'b0000000001000000: n9585_o = n9584_o;
      16'b0000000000100000: n9585_o = n9584_o;
      16'b0000000000010000: n9585_o = n9584_o;
      16'b0000000000001000: n9585_o = n9584_o;
      16'b0000000000000100: n9585_o = n9584_o;
      16'b0000000000000010: n9585_o = n9584_o;
      16'b0000000000000001: n9585_o = n9584_o;
      default: n9585_o = n9584_o;
    endcase
  assign n9586_o = sndopc[14];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9557_o)
      16'b1000000000000000: n9587_o = n9586_o;
      16'b0100000000000000: n9587_o = 1'b0;
      16'b0010000000000000: n9587_o = n9586_o;
      16'b0001000000000000: n9587_o = n9586_o;
      16'b0000100000000000: n9587_o = n9586_o;
      16'b0000010000000000: n9587_o = n9586_o;
      16'b0000001000000000: n9587_o = n9586_o;
      16'b0000000100000000: n9587_o = n9586_o;
      16'b0000000010000000: n9587_o = n9586_o;
      16'b0000000001000000: n9587_o = n9586_o;
      16'b0000000000100000: n9587_o = n9586_o;
      16'b0000000000010000: n9587_o = n9586_o;
      16'b0000000000001000: n9587_o = n9586_o;
      16'b0000000000000100: n9587_o = n9586_o;
      16'b0000000000000010: n9587_o = n9586_o;
      16'b0000000000000001: n9587_o = n9586_o;
      default: n9587_o = n9586_o;
    endcase
  assign n9588_o = sndopc[15];
  /* TG68KdotC_Kernel.vhd:4116:41  */
  always @*
    case (n9557_o)
      16'b1000000000000000: n9589_o = 1'b0;
      16'b0100000000000000: n9589_o = n9588_o;
      16'b0010000000000000: n9589_o = n9588_o;
      16'b0001000000000000: n9589_o = n9588_o;
      16'b0000100000000000: n9589_o = n9588_o;
      16'b0000010000000000: n9589_o = n9588_o;
      16'b0000001000000000: n9589_o = n9588_o;
      16'b0000000100000000: n9589_o = n9588_o;
      16'b0000000010000000: n9589_o = n9588_o;
      16'b0000000001000000: n9589_o = n9588_o;
      16'b0000000000100000: n9589_o = n9588_o;
      16'b0000000000010000: n9589_o = n9588_o;
      16'b0000000000001000: n9589_o = n9588_o;
      16'b0000000000000100: n9589_o = n9588_o;
      16'b0000000000000010: n9589_o = n9588_o;
      16'b0000000000000001: n9589_o = n9588_o;
      default: n9589_o = n9588_o;
    endcase
  assign n9590_o = {n9589_o, n9587_o, n9585_o, n9583_o, n9581_o, n9579_o, n9577_o, n9575_o, n9573_o, n9571_o, n9569_o, n9567_o, n9565_o, n9563_o, n9561_o, n9559_o};
  /* TG68KdotC_Kernel.vhd:4115:33  */
  assign n9591_o = n9508_o ? n9590_o : sndopc;
  /* TG68KdotC_Kernel.vhd:4113:33  */
  assign n9592_o = decodeopc ? n9505_o : n9591_o;
  /* TG68KdotC_Kernel.vhd:4144:26  */
  assign n9600_o = sndopc[3:0];
  /* TG68KdotC_Kernel.vhd:4144:38  */
  assign n9602_o = n9600_o == 4'b0000;
  /* TG68KdotC_Kernel.vhd:4145:34  */
  assign n9603_o = sndopc[7:4];
  /* TG68KdotC_Kernel.vhd:4145:46  */
  assign n9605_o = n9603_o == 4'b0000;
  /* TG68KdotC_Kernel.vhd:4147:42  */
  assign n9607_o = sndopc[11:8];
  /* TG68KdotC_Kernel.vhd:4147:55  */
  assign n9609_o = n9607_o == 4'b0000;
  /* TG68KdotC_Kernel.vhd:4148:50  */
  assign n9610_o = sndopc[15:12];
  /* TG68KdotC_Kernel.vhd:4148:64  */
  assign n9612_o = n9610_o == 4'b0000;
  /* TG68KdotC_Kernel.vhd:4148:41  */
  assign n9615_o = n9612_o ? 1'b0 : 1'b1;
  /* TG68KdotC_Kernel.vhd:4152:60  */
  assign n9617_o = sndopc[15:12];
  /* TG68KdotC_Kernel.vhd:4154:60  */
  assign n9618_o = sndopc[11:8];
  /* TG68KdotC_Kernel.vhd:4147:33  */
  assign n9620_o = n9609_o ? 1'b1 : 1'b0;
  /* TG68KdotC_Kernel.vhd:4147:33  */
  assign n9621_o = n9609_o ? n9617_o : n9618_o;
  /* TG68KdotC_Kernel.vhd:4147:33  */
  assign n9623_o = n9609_o ? n9615_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:4157:52  */
  assign n9624_o = sndopc[7:4];
  assign n9626_o = {1'b1, n9620_o};
  assign n9627_o = n9626_o[0];
  /* TG68KdotC_Kernel.vhd:4145:25  */
  assign n9628_o = n9605_o ? n9627_o : 1'b1;
  assign n9629_o = n9626_o[1];
  /* TG68KdotC_Kernel.vhd:4145:25  */
  assign n9631_o = n9605_o ? n9629_o : 1'b0;
  /* TG68KdotC_Kernel.vhd:4145:25  */
  assign n9632_o = n9605_o ? n9621_o : n9624_o;
  /* TG68KdotC_Kernel.vhd:4145:25  */
  assign n9634_o = n9605_o ? n9623_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:4161:44  */
  assign n9635_o = sndopc[3:0];
  assign n9636_o = {n9631_o, n9628_o};
  /* TG68KdotC_Kernel.vhd:4144:17  */
  assign n9638_o = n9602_o ? n9636_o : 2'b00;
  /* TG68KdotC_Kernel.vhd:4144:17  */
  assign n9641_o = n9602_o ? n9632_o : n9635_o;
  /* TG68KdotC_Kernel.vhd:4144:17  */
  assign n9643_o = n9602_o ? n9634_o : 1'b1;
  /* TG68KdotC_Kernel.vhd:4163:29  */
  assign n9645_o = movem_mux[1:0];
  /* TG68KdotC_Kernel.vhd:4163:41  */
  assign n9647_o = n9645_o == 2'b00;
  /* TG68KdotC_Kernel.vhd:4165:37  */
  assign n9649_o = movem_mux[2];
  /* TG68KdotC_Kernel.vhd:4165:40  */
  assign n9650_o = ~n9649_o;
  assign n9652_o = n9639_o[0];
  /* TG68KdotC_Kernel.vhd:4165:25  */
  assign n9653_o = n9650_o ? 1'b1 : n9652_o;
  /* TG68KdotC_Kernel.vhd:4169:37  */
  assign n9654_o = movem_mux[0];
  /* TG68KdotC_Kernel.vhd:4169:40  */
  assign n9655_o = ~n9654_o;
  assign n9657_o = n9639_o[0];
  /* TG68KdotC_Kernel.vhd:4169:25  */
  assign n9658_o = n9655_o ? 1'b1 : n9657_o;
  assign n9659_o = {1'b1, n9653_o};
  assign n9660_o = n9659_o[0];
  /* TG68KdotC_Kernel.vhd:4163:17  */
  assign n9661_o = n9647_o ? n9660_o : n9658_o;
  assign n9662_o = n9659_o[1];
  assign n9663_o = n9639_o[1];
  /* TG68KdotC_Kernel.vhd:4163:17  */
  assign n9664_o = n9647_o ? n9662_o : n9663_o;
  /* TG68KdotC_Kernel.vhd:464:17  */
  always @(posedge clk)
    n9667_q <= n125_o;
  /* TG68KdotC_Kernel.vhd:458:17  */
  assign n9668_o = clkena_in ? n106_o : syncreset;
  /* TG68KdotC_Kernel.vhd:458:17  */
  always @(posedge clk or posedge n102_o)
    if (n102_o)
      n9669_q <= 4'b0000;
    else
      n9669_q <= n9668_o;
  /* TG68KdotC_Kernel.vhd:458:17  */
  assign n9670_o = clkena_in ? n108_o : reset;
  /* TG68KdotC_Kernel.vhd:458:17  */
  always @(posedge clk or posedge n102_o)
    if (n102_o)
      n9671_q <= 1'b1;
    else
      n9671_q <= n9670_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9672_q <= n1512_o;
  /* TG68KdotC_Kernel.vhd:947:17  */
  assign n9673_o = n1062_o ? addr : tmp_tg68_pc;
  /* TG68KdotC_Kernel.vhd:947:17  */
  always @(posedge clk)
    n9674_q <= n9673_o;
  /* TG68KdotC_Kernel.vhd:947:17  */
  assign n9675_o = n1063_o ? addr : memaddr;
  /* TG68KdotC_Kernel.vhd:947:17  */
  always @(posedge clk)
    n9676_q <= n9675_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9677_q <= n1514_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9678_q <= n1515_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9679_q <= n1517_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9680_q <= n1519_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9681_q <= n1520_o;
  /* TG68KdotC_Kernel.vhd:4110:17  */
  assign n9682_o = clkena_lw ? n9592_o : sndopc;
  /* TG68KdotC_Kernel.vhd:4110:17  */
  always @(posedge clk)
    n9683_q <= n9682_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9684_q <= n1521_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9685_q <= n1522_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9686_q <= n1524_o;
  /* TG68KdotC_Kernel.vhd:560:17  */
  assign n9688_o = clkena_lw ? rf_source_addr : rf_source_addrd;
  /* TG68KdotC_Kernel.vhd:560:17  */
  always @(posedge clk)
    n9689_q <= n9688_o;
  /* TG68KdotC_Kernel.vhd:560:17  */
  assign n9690_o = {n356_o, n335_o, n353_o};
  /* TG68KdotC_Kernel.vhd:560:17  */
  assign n9693_o = clkena_lw ? rf_dest_addr : rdindex_a;
  /* TG68KdotC_Kernel.vhd:560:17  */
  always @(posedge clk)
    n9694_q <= n9693_o;
  /* TG68KdotC_Kernel.vhd:560:17  */
  assign n9695_o = clkena_lw ? rf_source_addr : rdindex_b;
  /* TG68KdotC_Kernel.vhd:560:17  */
  always @(posedge clk)
    n9696_q <= n9695_o;
  /* TG68KdotC_Kernel.vhd:560:17  */
  assign n9697_o = clkena_lw ? n291_o : wr_areg;
  /* TG68KdotC_Kernel.vhd:560:17  */
  always @(posedge clk)
    n9698_q <= n9697_o;
  /* TG68KdotC_Kernel.vhd:947:17  */
  assign n9699_o = clkena_in ? n1049_o : memaddr_delta_rega;
  /* TG68KdotC_Kernel.vhd:947:17  */
  always @(posedge clk)
    n9700_q <= n9699_o;
  /* TG68KdotC_Kernel.vhd:947:17  */
  assign n9701_o = clkena_in ? n1051_o : memaddr_delta_regb;
  /* TG68KdotC_Kernel.vhd:947:17  */
  always @(posedge clk)
    n9702_q <= n9701_o;
  /* TG68KdotC_Kernel.vhd:947:17  */
  assign n9703_o = clkena_in ? n1054_o : use_base;
  /* TG68KdotC_Kernel.vhd:947:17  */
  always @(posedge clk)
    n9704_q <= n9703_o;
  /* TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9705_q <= n790_o;
  /* TG68KdotC_Kernel.vhd:743:9  */
  assign n9706_o = {n619_o, n626_o};
  /* TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9708_q <= n791_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9709_q <= n1525_o;
  assign n9711_o = {n987_o, n984_o};
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9712_q <= n1527_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9713_q <= n1528_o;
  /* TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9714_q <= n793_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9715_q <= n1530_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9716_q <= n1532_o;
  /* TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9717_q <= n795_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9718_q <= n1534_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9719_q <= n1536_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9720_q <= n1538_o;
  /* TG68KdotC_Kernel.vhd:1370:17  */
  always @(posedge clk)
    n9721_q <= n1884_o;
  /* TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9722_q <= n796_o;
  /* TG68KdotC_Kernel.vhd:1260:17  */
  assign n9723_o = clkena_lw ? n1647_o : exec_tas;
  /* TG68KdotC_Kernel.vhd:1260:17  */
  always @(posedge clk)
    n9724_q <= n9723_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9725_q <= n1539_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9726_q <= n1541_o;
  /* TG68KdotC_Kernel.vhd:4110:17  */
  assign n9727_o = clkena_lw ? n9504_o : movem_actiond;
  /* TG68KdotC_Kernel.vhd:4110:17  */
  always @(posedge clk)
    n9728_q <= n9727_o;
  /* TG68KdotC_Kernel.vhd:4110:17  */
  assign n9729_o = {n9638_o, n9664_o, n9661_o};
  /* TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9731_q <= n798_o;
  /* TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9732_q <= n800_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9733_q <= n1543_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9734_q <= n1545_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9735_q <= n1547_o;
  /* TG68KdotC_Kernel.vhd:3254:17  */
  always @(posedge clk)
    n9736_q <= n8007_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9737_q <= n1548_o;
  /* TG68KdotC_Kernel.vhd:1370:17  */
  always @(posedge clk)
    n9738_q <= n1886_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9739_q <= n1550_o;
  /* TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9740_q <= n801_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9741_q <= n1552_o;
  /* TG68KdotC_Kernel.vhd:876:17  */
  assign n9742_o = clkena_lw ? n913_o : trap_vector;
  /* TG68KdotC_Kernel.vhd:876:17  */
  always @(posedge clk)
    n9743_q <= n9742_o;
  /* TG68KdotC_Kernel.vhd:560:17  */
  assign n9744_o = n306_o ? reg_qa : usp;
  /* TG68KdotC_Kernel.vhd:560:17  */
  always @(posedge clk)
    n9745_q <= n9744_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9746_q <= n1553_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9747_q <= n1554_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9748_q <= n1556_o;
  /* TG68KdotC_Kernel.vhd:1370:17  */
  always @(posedge clk)
    n9749_q <= n1888_o;
  /* TG68KdotC_Kernel.vhd:1370:17  */
  always @(posedge clk)
    n9750_q <= n1890_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9751_q <= n1558_o;
  /* TG68KdotC_Kernel.vhd:743:9  */
  always @(posedge clk)
    n9752_q <= n803_o;
  /* TG68KdotC_Kernel.vhd:743:9  */
  assign n9753_o = {n169_o, n172_o};
  /* TG68KdotC_Kernel.vhd:484:17  */
  assign n9754_o = n176_o ? n181_o : bf_ext_in;
  /* TG68KdotC_Kernel.vhd:484:17  */
  always @(posedge clk)
    n9755_q <= n9754_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9756_q <= n1560_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9757_q <= n1561_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9758_q <= n1562_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9759_q <= n1563_o;
  /* TG68KdotC_Kernel.vhd:1260:17  */
  always @(posedge clk)
    n9760_q <= n1617_o;
  /* TG68KdotC_Kernel.vhd:484:17  */
  always @(posedge clk)
    n9761_q <= n228_o;
  /* TG68KdotC_Kernel.vhd:484:17  */
  always @(posedge clk)
    n9762_q <= n229_o;
  /* TG68KdotC_Kernel.vhd:484:17  */
  assign n9763_o = {n1744_o, n1741_o, n1747_o};
  assign n9764_o = {1'b0, n1691_o};
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9765_q <= n1564_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9766_q <= n1565_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  assign n9767_o = {1'b0, n1704_o};
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9768_q <= n1566_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9769_q <= n1567_o;
  /* TG68KdotC_Kernel.vhd:4045:9  */
  always @(posedge clk)
    n9770_q <= n9366_o;
  /* TG68KdotC_Kernel.vhd:4045:9  */
  always @(posedge clk)
    n9771_q <= n9368_o;
  /* TG68KdotC_Kernel.vhd:4045:9  */
  always @(posedge clk)
    n9772_q <= n9369_o;
  /* TG68KdotC_Kernel.vhd:4045:9  */
  always @(posedge clk)
    n9773_q <= n9370_o;
  /* TG68KdotC_Kernel.vhd:4045:9  */
  assign n9774_o = {n9235_o, n9233_o, n9231_o, n9227_o, n9223_o, n9219_o, n9218_o, n7836_o, n7813_o, n9217_o, n9272_o, n9271_o, n9215_o, n9211_o, n7808_o, n9210_o, n9209_o, n9208_o, n9206_o, n9264_o, n9204_o, n9267_o, n9200_o, n9261_o, n9199_o, n9195_o, n9191_o, n9187_o, n9252_o, n9183_o, n9182_o, n9246_o, n9178_o, n9177_o, n9176_o, n7800_o, n2002_o, n9175_o, n9171_o, n9167_o, n9166_o, n9240_o, n9162_o, n9161_o, n7826_o, n7793_o, n9237_o, n9160_o, n9158_o, n9157_o, n9156_o, n7821_o, n9155_o, n9154_o, n9152_o, n7787_o, n7820_o, n9150_o};
  assign n9775_o = {n7852_o, n7863_o, n7850_o, n7862_o, n7996_o, n7906_o, n7860_o, n7995_o, n7858_o, n7994_o, n9282_o, n9281_o, n9283_o, n7842_o};
  /* TG68KdotC_Kernel.vhd:1260:17  */
  assign n9776_o = clkena_lw ? n1661_o : exec;
  /* TG68KdotC_Kernel.vhd:1260:17  */
  always @(posedge clk)
    n9777_q <= n9776_o;
  /* TG68KdotC_Kernel.vhd:3254:17  */
  always @(posedge clk)
    n9778_q <= n8009_o;
  /* TG68KdotC_Kernel.vhd:1370:17  */
  always @(posedge clk)
    n9779_q <= n1882_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  always @(posedge clk)
    n9780_q <= n1510_o;
  /* TG68KdotC_Kernel.vhd:1059:17  */
  assign n9781_o = {n9779_q, n9780_q};
  /* TG68KdotC_Kernel.vhd:558:35  */
  reg [31:0] regfile[15:0] ; // memory
  initial begin
    regfile[15] = 32'b00000000000000000000000000000000;
    regfile[14] = 32'b00000000000000000000000000000000;
    regfile[13] = 32'b00000000000000000000000000000000;
    regfile[12] = 32'b00000000000000000000000000000000;
    regfile[11] = 32'b00000000000000000000000000000000;
    regfile[10] = 32'b00000000000000000000000000000000;
    regfile[9] = 32'b00000000000000000000000000000000;
    regfile[8] = 32'b00000000000000000000000000000000;
    regfile[7] = 32'b00000000000000000000000000000000;
    regfile[6] = 32'b00000000000000000000000000000000;
    regfile[5] = 32'b00000000000000000000000000000000;
    regfile[4] = 32'b00000000000000000000000000000000;
    regfile[3] = 32'b00000000000000000000000000000000;
    regfile[2] = 32'b00000000000000000000000000000000;
    regfile[1] = 32'b00000000000000000000000000000000;
    regfile[0] = 32'b00000000000000000000000000000000;
    end
  assign n9783_data = regfile[rdindex_b];
  assign n9784_data = regfile[rdindex_a];
  always @(posedge clk)
    if (n302_o)
      regfile[rdindex_a] <= regin;
  /* TG68KdotC_Kernel.vhd:559:35  */
  /* TG68KdotC_Kernel.vhd:558:35  */
  /* TG68KdotC_Kernel.vhd:567:49  */
endmodule

module tg68kdotc_verilog_wrapper
  (input  clk,
   input  nReset,
   input  clkena_in,
   input  [15:0] data_in,
   input  [2:0] IPL,
   input  IPL_autovector,
   input  berr,
   output [31:0] addr_out,
   output [2:0] FC,
   output [15:0] data_write,
   output [1:0] busstate,
   output nWr,
   output nUDS,
   output nLDS,
   output nResetOut,
   output skipFetch);
  wire [31:0] tg68kdotcinst_addr_out;
  wire [15:0] tg68kdotcinst_data_write;
  wire tg68kdotcinst_nwr;
  wire tg68kdotcinst_nuds;
  wire tg68kdotcinst_nlds;
  wire [1:0] tg68kdotcinst_busstate;
  wire tg68kdotcinst_longword;
  wire tg68kdotcinst_nresetout;
  wire [2:0] tg68kdotcinst_fc;
  wire tg68kdotcinst_clr_berr;
  wire tg68kdotcinst_skipfetch;
  wire [31:0] tg68kdotcinst_regin_out;
  wire [3:0] tg68kdotcinst_cacr_out;
  wire [31:0] tg68kdotcinst_vbr_out;
  localparam [1:0] n9_o = 2'b01;
  assign addr_out = tg68kdotcinst_addr_out;
  assign FC = tg68kdotcinst_fc;
  assign data_write = tg68kdotcinst_data_write;
  assign busstate = tg68kdotcinst_busstate;
  assign nWr = tg68kdotcinst_nwr;
  assign nUDS = tg68kdotcinst_nuds;
  assign nLDS = tg68kdotcinst_nlds;
  assign nResetOut = tg68kdotcinst_nresetout;
  assign skipFetch = tg68kdotcinst_skipfetch;
  /* tg68dotc_verilog_wrapper.vhd:27:3  */
  tg68kdotc_kernel_0_2_2_2_2_2_0_0 tg68kdotcinst (
    .clk(clk),
    .nreset(nReset),
    .clkena_in(clkena_in),
    .data_in(data_in),
    .ipl(IPL),
    .ipl_autovector(IPL_autovector),
    .berr(berr),
    .cpu(n9_o),
    .addr_out(tg68kdotcinst_addr_out),
    .data_write(tg68kdotcinst_data_write),
    .nwr(tg68kdotcinst_nwr),
    .nuds(tg68kdotcinst_nuds),
    .nlds(tg68kdotcinst_nlds),
    .busstate(tg68kdotcinst_busstate),
    .longword(),
    .nresetout(tg68kdotcinst_nresetout),
    .fc(tg68kdotcinst_fc),
    .clr_berr(),
    .skipfetch(tg68kdotcinst_skipfetch),
    .regin_out(),
    .cacr_out(),
    .vbr_out());
endmodule

