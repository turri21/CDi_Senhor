
function signed [17:0] PLM_AUDIO_SYNTHESIS_WINDOW(bit [8:0] index);
    case (index)
        0:   PLM_AUDIO_SYNTHESIS_WINDOW = 0;
        1:   PLM_AUDIO_SYNTHESIS_WINDOW = -1;
        2:   PLM_AUDIO_SYNTHESIS_WINDOW = -1;
        3:   PLM_AUDIO_SYNTHESIS_WINDOW = -1;
        4:   PLM_AUDIO_SYNTHESIS_WINDOW = -1;
        5:   PLM_AUDIO_SYNTHESIS_WINDOW = -1;
        6:   PLM_AUDIO_SYNTHESIS_WINDOW = -1;
        7:   PLM_AUDIO_SYNTHESIS_WINDOW = -2;
        8:   PLM_AUDIO_SYNTHESIS_WINDOW = -2;
        9:   PLM_AUDIO_SYNTHESIS_WINDOW = -2;
        10:  PLM_AUDIO_SYNTHESIS_WINDOW = -2;
        11:  PLM_AUDIO_SYNTHESIS_WINDOW = -3;
        12:  PLM_AUDIO_SYNTHESIS_WINDOW = -3;
        13:  PLM_AUDIO_SYNTHESIS_WINDOW = -4;
        14:  PLM_AUDIO_SYNTHESIS_WINDOW = -4;
        15:  PLM_AUDIO_SYNTHESIS_WINDOW = -5;
        16:  PLM_AUDIO_SYNTHESIS_WINDOW = -5;
        17:  PLM_AUDIO_SYNTHESIS_WINDOW = -6;
        18:  PLM_AUDIO_SYNTHESIS_WINDOW = -7;
        19:  PLM_AUDIO_SYNTHESIS_WINDOW = -7;
        20:  PLM_AUDIO_SYNTHESIS_WINDOW = -8;
        21:  PLM_AUDIO_SYNTHESIS_WINDOW = -9;
        22:  PLM_AUDIO_SYNTHESIS_WINDOW = -10;
        23:  PLM_AUDIO_SYNTHESIS_WINDOW = -11;
        24:  PLM_AUDIO_SYNTHESIS_WINDOW = -13;
        25:  PLM_AUDIO_SYNTHESIS_WINDOW = -14;
        26:  PLM_AUDIO_SYNTHESIS_WINDOW = -16;
        27:  PLM_AUDIO_SYNTHESIS_WINDOW = -17;
        28:  PLM_AUDIO_SYNTHESIS_WINDOW = -19;
        29:  PLM_AUDIO_SYNTHESIS_WINDOW = -21;
        30:  PLM_AUDIO_SYNTHESIS_WINDOW = -24;
        31:  PLM_AUDIO_SYNTHESIS_WINDOW = -26;
        32:  PLM_AUDIO_SYNTHESIS_WINDOW = -29;
        33:  PLM_AUDIO_SYNTHESIS_WINDOW = -31;
        34:  PLM_AUDIO_SYNTHESIS_WINDOW = -35;
        35:  PLM_AUDIO_SYNTHESIS_WINDOW = -38;
        36:  PLM_AUDIO_SYNTHESIS_WINDOW = -41;
        37:  PLM_AUDIO_SYNTHESIS_WINDOW = -45;
        38:  PLM_AUDIO_SYNTHESIS_WINDOW = -49;
        39:  PLM_AUDIO_SYNTHESIS_WINDOW = -53;
        40:  PLM_AUDIO_SYNTHESIS_WINDOW = -58;
        41:  PLM_AUDIO_SYNTHESIS_WINDOW = -63;
        42:  PLM_AUDIO_SYNTHESIS_WINDOW = -68;
        43:  PLM_AUDIO_SYNTHESIS_WINDOW = -73;
        44:  PLM_AUDIO_SYNTHESIS_WINDOW = -79;
        45:  PLM_AUDIO_SYNTHESIS_WINDOW = -85;
        46:  PLM_AUDIO_SYNTHESIS_WINDOW = -91;
        47:  PLM_AUDIO_SYNTHESIS_WINDOW = -97;
        48:  PLM_AUDIO_SYNTHESIS_WINDOW = -104;
        49:  PLM_AUDIO_SYNTHESIS_WINDOW = -111;
        50:  PLM_AUDIO_SYNTHESIS_WINDOW = -117;
        51:  PLM_AUDIO_SYNTHESIS_WINDOW = -125;
        52:  PLM_AUDIO_SYNTHESIS_WINDOW = -132;
        53:  PLM_AUDIO_SYNTHESIS_WINDOW = -139;
        54:  PLM_AUDIO_SYNTHESIS_WINDOW = -147;
        55:  PLM_AUDIO_SYNTHESIS_WINDOW = -154;
        56:  PLM_AUDIO_SYNTHESIS_WINDOW = -161;
        57:  PLM_AUDIO_SYNTHESIS_WINDOW = -169;
        58:  PLM_AUDIO_SYNTHESIS_WINDOW = -176;
        59:  PLM_AUDIO_SYNTHESIS_WINDOW = -183;
        60:  PLM_AUDIO_SYNTHESIS_WINDOW = -190;
        61:  PLM_AUDIO_SYNTHESIS_WINDOW = -196;
        62:  PLM_AUDIO_SYNTHESIS_WINDOW = -202;
        63:  PLM_AUDIO_SYNTHESIS_WINDOW = -208;
        64:  PLM_AUDIO_SYNTHESIS_WINDOW = 213;
        65:  PLM_AUDIO_SYNTHESIS_WINDOW = 218;
        66:  PLM_AUDIO_SYNTHESIS_WINDOW = 222;
        67:  PLM_AUDIO_SYNTHESIS_WINDOW = 225;
        68:  PLM_AUDIO_SYNTHESIS_WINDOW = 227;
        69:  PLM_AUDIO_SYNTHESIS_WINDOW = 228;
        70:  PLM_AUDIO_SYNTHESIS_WINDOW = 228;
        71:  PLM_AUDIO_SYNTHESIS_WINDOW = 227;
        72:  PLM_AUDIO_SYNTHESIS_WINDOW = 224;
        73:  PLM_AUDIO_SYNTHESIS_WINDOW = 221;
        74:  PLM_AUDIO_SYNTHESIS_WINDOW = 215;
        75:  PLM_AUDIO_SYNTHESIS_WINDOW = 208;
        76:  PLM_AUDIO_SYNTHESIS_WINDOW = 200;
        77:  PLM_AUDIO_SYNTHESIS_WINDOW = 189;
        78:  PLM_AUDIO_SYNTHESIS_WINDOW = 177;
        79:  PLM_AUDIO_SYNTHESIS_WINDOW = 163;
        80:  PLM_AUDIO_SYNTHESIS_WINDOW = 146;
        81:  PLM_AUDIO_SYNTHESIS_WINDOW = 127;
        82:  PLM_AUDIO_SYNTHESIS_WINDOW = 106;
        83:  PLM_AUDIO_SYNTHESIS_WINDOW = 83;
        84:  PLM_AUDIO_SYNTHESIS_WINDOW = 57;
        85:  PLM_AUDIO_SYNTHESIS_WINDOW = 29;
        86:  PLM_AUDIO_SYNTHESIS_WINDOW = -2;
        87:  PLM_AUDIO_SYNTHESIS_WINDOW = -36;
        88:  PLM_AUDIO_SYNTHESIS_WINDOW = -72;
        89:  PLM_AUDIO_SYNTHESIS_WINDOW = -111;
        90:  PLM_AUDIO_SYNTHESIS_WINDOW = -153;
        91:  PLM_AUDIO_SYNTHESIS_WINDOW = -197;
        92:  PLM_AUDIO_SYNTHESIS_WINDOW = -244;
        93:  PLM_AUDIO_SYNTHESIS_WINDOW = -294;
        94:  PLM_AUDIO_SYNTHESIS_WINDOW = -347;
        95:  PLM_AUDIO_SYNTHESIS_WINDOW = -401;
        96:  PLM_AUDIO_SYNTHESIS_WINDOW = -459;
        97:  PLM_AUDIO_SYNTHESIS_WINDOW = -519;
        98:  PLM_AUDIO_SYNTHESIS_WINDOW = -581;
        99:  PLM_AUDIO_SYNTHESIS_WINDOW = -645;
        100: PLM_AUDIO_SYNTHESIS_WINDOW = -711;
        101: PLM_AUDIO_SYNTHESIS_WINDOW = -779;
        102: PLM_AUDIO_SYNTHESIS_WINDOW = -848;
        103: PLM_AUDIO_SYNTHESIS_WINDOW = -919;
        104: PLM_AUDIO_SYNTHESIS_WINDOW = -991;
        105: PLM_AUDIO_SYNTHESIS_WINDOW = -1064;
        106: PLM_AUDIO_SYNTHESIS_WINDOW = -1137;
        107: PLM_AUDIO_SYNTHESIS_WINDOW = -1210;
        108: PLM_AUDIO_SYNTHESIS_WINDOW = -1283;
        109: PLM_AUDIO_SYNTHESIS_WINDOW = -1356;
        110: PLM_AUDIO_SYNTHESIS_WINDOW = -1428;
        111: PLM_AUDIO_SYNTHESIS_WINDOW = -1498;
        112: PLM_AUDIO_SYNTHESIS_WINDOW = -1567;
        113: PLM_AUDIO_SYNTHESIS_WINDOW = -1634;
        114: PLM_AUDIO_SYNTHESIS_WINDOW = -1698;
        115: PLM_AUDIO_SYNTHESIS_WINDOW = -1759;
        116: PLM_AUDIO_SYNTHESIS_WINDOW = -1817;
        117: PLM_AUDIO_SYNTHESIS_WINDOW = -1870;
        118: PLM_AUDIO_SYNTHESIS_WINDOW = -1919;
        119: PLM_AUDIO_SYNTHESIS_WINDOW = -1962;
        120: PLM_AUDIO_SYNTHESIS_WINDOW = -2001;
        121: PLM_AUDIO_SYNTHESIS_WINDOW = -2032;
        122: PLM_AUDIO_SYNTHESIS_WINDOW = -2057;
        123: PLM_AUDIO_SYNTHESIS_WINDOW = -2075;
        124: PLM_AUDIO_SYNTHESIS_WINDOW = -2085;
        125: PLM_AUDIO_SYNTHESIS_WINDOW = -2087;
        126: PLM_AUDIO_SYNTHESIS_WINDOW = -2080;
        127: PLM_AUDIO_SYNTHESIS_WINDOW = -2063;
        128: PLM_AUDIO_SYNTHESIS_WINDOW = 2037;
        129: PLM_AUDIO_SYNTHESIS_WINDOW = 2000;
        130: PLM_AUDIO_SYNTHESIS_WINDOW = 1952;
        131: PLM_AUDIO_SYNTHESIS_WINDOW = 1893;
        132: PLM_AUDIO_SYNTHESIS_WINDOW = 1822;
        133: PLM_AUDIO_SYNTHESIS_WINDOW = 1739;
        134: PLM_AUDIO_SYNTHESIS_WINDOW = 1644;
        135: PLM_AUDIO_SYNTHESIS_WINDOW = 1535;
        136: PLM_AUDIO_SYNTHESIS_WINDOW = 1414;
        137: PLM_AUDIO_SYNTHESIS_WINDOW = 1280;
        138: PLM_AUDIO_SYNTHESIS_WINDOW = 1131;
        139: PLM_AUDIO_SYNTHESIS_WINDOW = 970;
        140: PLM_AUDIO_SYNTHESIS_WINDOW = 794;
        141: PLM_AUDIO_SYNTHESIS_WINDOW = 605;
        142: PLM_AUDIO_SYNTHESIS_WINDOW = 402;
        143: PLM_AUDIO_SYNTHESIS_WINDOW = 185;
        144: PLM_AUDIO_SYNTHESIS_WINDOW = -45;
        145: PLM_AUDIO_SYNTHESIS_WINDOW = -288;
        146: PLM_AUDIO_SYNTHESIS_WINDOW = -545;
        147: PLM_AUDIO_SYNTHESIS_WINDOW = -814;
        148: PLM_AUDIO_SYNTHESIS_WINDOW = -1095;
        149: PLM_AUDIO_SYNTHESIS_WINDOW = -1388;
        150: PLM_AUDIO_SYNTHESIS_WINDOW = -1692;
        151: PLM_AUDIO_SYNTHESIS_WINDOW = -2006;
        152: PLM_AUDIO_SYNTHESIS_WINDOW = -2330;
        153: PLM_AUDIO_SYNTHESIS_WINDOW = -2663;
        154: PLM_AUDIO_SYNTHESIS_WINDOW = -3004;
        155: PLM_AUDIO_SYNTHESIS_WINDOW = -3351;
        156: PLM_AUDIO_SYNTHESIS_WINDOW = -3705;
        157: PLM_AUDIO_SYNTHESIS_WINDOW = -4063;
        158: PLM_AUDIO_SYNTHESIS_WINDOW = -4425;
        159: PLM_AUDIO_SYNTHESIS_WINDOW = -4788;
        160: PLM_AUDIO_SYNTHESIS_WINDOW = -5153;
        161: PLM_AUDIO_SYNTHESIS_WINDOW = -5517;
        162: PLM_AUDIO_SYNTHESIS_WINDOW = -5879;
        163: PLM_AUDIO_SYNTHESIS_WINDOW = -6237;
        164: PLM_AUDIO_SYNTHESIS_WINDOW = -6589;
        165: PLM_AUDIO_SYNTHESIS_WINDOW = -6935;
        166: PLM_AUDIO_SYNTHESIS_WINDOW = -7271;
        167: PLM_AUDIO_SYNTHESIS_WINDOW = -7597;
        168: PLM_AUDIO_SYNTHESIS_WINDOW = -7910;
        169: PLM_AUDIO_SYNTHESIS_WINDOW = -8209;
        170: PLM_AUDIO_SYNTHESIS_WINDOW = -8491;
        171: PLM_AUDIO_SYNTHESIS_WINDOW = -8755;
        172: PLM_AUDIO_SYNTHESIS_WINDOW = -8998;
        173: PLM_AUDIO_SYNTHESIS_WINDOW = -9219;
        174: PLM_AUDIO_SYNTHESIS_WINDOW = -9416;
        175: PLM_AUDIO_SYNTHESIS_WINDOW = -9585;
        176: PLM_AUDIO_SYNTHESIS_WINDOW = -9727;
        177: PLM_AUDIO_SYNTHESIS_WINDOW = -9838;
        178: PLM_AUDIO_SYNTHESIS_WINDOW = -9916;
        179: PLM_AUDIO_SYNTHESIS_WINDOW = -9959;
        180: PLM_AUDIO_SYNTHESIS_WINDOW = -9966;
        181: PLM_AUDIO_SYNTHESIS_WINDOW = -9935;
        182: PLM_AUDIO_SYNTHESIS_WINDOW = -9863;
        183: PLM_AUDIO_SYNTHESIS_WINDOW = -9750;
        184: PLM_AUDIO_SYNTHESIS_WINDOW = -9592;
        185: PLM_AUDIO_SYNTHESIS_WINDOW = -9389;
        186: PLM_AUDIO_SYNTHESIS_WINDOW = -9139;
        187: PLM_AUDIO_SYNTHESIS_WINDOW = -8840;
        188: PLM_AUDIO_SYNTHESIS_WINDOW = -8492;
        189: PLM_AUDIO_SYNTHESIS_WINDOW = -8092;
        190: PLM_AUDIO_SYNTHESIS_WINDOW = -7640;
        191: PLM_AUDIO_SYNTHESIS_WINDOW = -7134;
        192: PLM_AUDIO_SYNTHESIS_WINDOW = 6574;
        193: PLM_AUDIO_SYNTHESIS_WINDOW = 5959;
        194: PLM_AUDIO_SYNTHESIS_WINDOW = 5288;
        195: PLM_AUDIO_SYNTHESIS_WINDOW = 4561;
        196: PLM_AUDIO_SYNTHESIS_WINDOW = 3776;
        197: PLM_AUDIO_SYNTHESIS_WINDOW = 2935;
        198: PLM_AUDIO_SYNTHESIS_WINDOW = 2037;
        199: PLM_AUDIO_SYNTHESIS_WINDOW = 1082;
        200: PLM_AUDIO_SYNTHESIS_WINDOW = 70;
        201: PLM_AUDIO_SYNTHESIS_WINDOW = -998;
        202: PLM_AUDIO_SYNTHESIS_WINDOW = -2122;
        203: PLM_AUDIO_SYNTHESIS_WINDOW = -3300;
        204: PLM_AUDIO_SYNTHESIS_WINDOW = -4533;
        205: PLM_AUDIO_SYNTHESIS_WINDOW = -5818;
        206: PLM_AUDIO_SYNTHESIS_WINDOW = -7154;
        207: PLM_AUDIO_SYNTHESIS_WINDOW = -8540;
        208: PLM_AUDIO_SYNTHESIS_WINDOW = -9975;
        209: PLM_AUDIO_SYNTHESIS_WINDOW = -11455;
        210: PLM_AUDIO_SYNTHESIS_WINDOW = -12980;
        211: PLM_AUDIO_SYNTHESIS_WINDOW = -14548;
        212: PLM_AUDIO_SYNTHESIS_WINDOW = -16155;
        213: PLM_AUDIO_SYNTHESIS_WINDOW = -17799;
        214: PLM_AUDIO_SYNTHESIS_WINDOW = -19478;
        215: PLM_AUDIO_SYNTHESIS_WINDOW = -21189;
        216: PLM_AUDIO_SYNTHESIS_WINDOW = -22929;
        217: PLM_AUDIO_SYNTHESIS_WINDOW = -24694;
        218: PLM_AUDIO_SYNTHESIS_WINDOW = -26482;
        219: PLM_AUDIO_SYNTHESIS_WINDOW = -28289;
        220: PLM_AUDIO_SYNTHESIS_WINDOW = -30112;
        221: PLM_AUDIO_SYNTHESIS_WINDOW = -31947;
        222: PLM_AUDIO_SYNTHESIS_WINDOW = -33791;
        223: PLM_AUDIO_SYNTHESIS_WINDOW = -35640;
        224: PLM_AUDIO_SYNTHESIS_WINDOW = -37489;
        225: PLM_AUDIO_SYNTHESIS_WINDOW = -39336;
        226: PLM_AUDIO_SYNTHESIS_WINDOW = -41176;
        227: PLM_AUDIO_SYNTHESIS_WINDOW = -43006;
        228: PLM_AUDIO_SYNTHESIS_WINDOW = -44821;
        229: PLM_AUDIO_SYNTHESIS_WINDOW = -46617;
        230: PLM_AUDIO_SYNTHESIS_WINDOW = -48390;
        231: PLM_AUDIO_SYNTHESIS_WINDOW = -50137;
        232: PLM_AUDIO_SYNTHESIS_WINDOW = -51853;
        233: PLM_AUDIO_SYNTHESIS_WINDOW = -53534;
        234: PLM_AUDIO_SYNTHESIS_WINDOW = -55178;
        235: PLM_AUDIO_SYNTHESIS_WINDOW = -56778;
        236: PLM_AUDIO_SYNTHESIS_WINDOW = -58333;
        237: PLM_AUDIO_SYNTHESIS_WINDOW = -59838;
        238: PLM_AUDIO_SYNTHESIS_WINDOW = -61289;
        239: PLM_AUDIO_SYNTHESIS_WINDOW = -62684;
        240: PLM_AUDIO_SYNTHESIS_WINDOW = -64019;
        241: PLM_AUDIO_SYNTHESIS_WINDOW = -65290;
        242: PLM_AUDIO_SYNTHESIS_WINDOW = -66494;
        243: PLM_AUDIO_SYNTHESIS_WINDOW = -67629;
        244: PLM_AUDIO_SYNTHESIS_WINDOW = -68692;
        245: PLM_AUDIO_SYNTHESIS_WINDOW = -69679;
        246: PLM_AUDIO_SYNTHESIS_WINDOW = -70590;
        247: PLM_AUDIO_SYNTHESIS_WINDOW = -71420;
        248: PLM_AUDIO_SYNTHESIS_WINDOW = -72169;
        249: PLM_AUDIO_SYNTHESIS_WINDOW = -72835;
        250: PLM_AUDIO_SYNTHESIS_WINDOW = -73415;
        251: PLM_AUDIO_SYNTHESIS_WINDOW = -73908;
        252: PLM_AUDIO_SYNTHESIS_WINDOW = -74313;
        253: PLM_AUDIO_SYNTHESIS_WINDOW = -74630;
        254: PLM_AUDIO_SYNTHESIS_WINDOW = -74856;
        255: PLM_AUDIO_SYNTHESIS_WINDOW = -74992;
        256: PLM_AUDIO_SYNTHESIS_WINDOW = 75038;
        257: PLM_AUDIO_SYNTHESIS_WINDOW = 74992;
        258: PLM_AUDIO_SYNTHESIS_WINDOW = 74856;
        259: PLM_AUDIO_SYNTHESIS_WINDOW = 74630;
        260: PLM_AUDIO_SYNTHESIS_WINDOW = 74313;
        261: PLM_AUDIO_SYNTHESIS_WINDOW = 73908;
        262: PLM_AUDIO_SYNTHESIS_WINDOW = 73415;
        263: PLM_AUDIO_SYNTHESIS_WINDOW = 72835;
        264: PLM_AUDIO_SYNTHESIS_WINDOW = 72169;
        265: PLM_AUDIO_SYNTHESIS_WINDOW = 71420;
        266: PLM_AUDIO_SYNTHESIS_WINDOW = 70590;
        267: PLM_AUDIO_SYNTHESIS_WINDOW = 69679;
        268: PLM_AUDIO_SYNTHESIS_WINDOW = 68692;
        269: PLM_AUDIO_SYNTHESIS_WINDOW = 67629;
        270: PLM_AUDIO_SYNTHESIS_WINDOW = 66494;
        271: PLM_AUDIO_SYNTHESIS_WINDOW = 65290;
        272: PLM_AUDIO_SYNTHESIS_WINDOW = 64019;
        273: PLM_AUDIO_SYNTHESIS_WINDOW = 62684;
        274: PLM_AUDIO_SYNTHESIS_WINDOW = 61289;
        275: PLM_AUDIO_SYNTHESIS_WINDOW = 59838;
        276: PLM_AUDIO_SYNTHESIS_WINDOW = 58333;
        277: PLM_AUDIO_SYNTHESIS_WINDOW = 56778;
        278: PLM_AUDIO_SYNTHESIS_WINDOW = 55178;
        279: PLM_AUDIO_SYNTHESIS_WINDOW = 53534;
        280: PLM_AUDIO_SYNTHESIS_WINDOW = 51853;
        281: PLM_AUDIO_SYNTHESIS_WINDOW = 50137;
        282: PLM_AUDIO_SYNTHESIS_WINDOW = 48390;
        283: PLM_AUDIO_SYNTHESIS_WINDOW = 46617;
        284: PLM_AUDIO_SYNTHESIS_WINDOW = 44821;
        285: PLM_AUDIO_SYNTHESIS_WINDOW = 43006;
        286: PLM_AUDIO_SYNTHESIS_WINDOW = 41176;
        287: PLM_AUDIO_SYNTHESIS_WINDOW = 39336;
        288: PLM_AUDIO_SYNTHESIS_WINDOW = 37489;
        289: PLM_AUDIO_SYNTHESIS_WINDOW = 35640;
        290: PLM_AUDIO_SYNTHESIS_WINDOW = 33791;
        291: PLM_AUDIO_SYNTHESIS_WINDOW = 31947;
        292: PLM_AUDIO_SYNTHESIS_WINDOW = 30112;
        293: PLM_AUDIO_SYNTHESIS_WINDOW = 28289;
        294: PLM_AUDIO_SYNTHESIS_WINDOW = 26482;
        295: PLM_AUDIO_SYNTHESIS_WINDOW = 24694;
        296: PLM_AUDIO_SYNTHESIS_WINDOW = 22929;
        297: PLM_AUDIO_SYNTHESIS_WINDOW = 21189;
        298: PLM_AUDIO_SYNTHESIS_WINDOW = 19478;
        299: PLM_AUDIO_SYNTHESIS_WINDOW = 17799;
        300: PLM_AUDIO_SYNTHESIS_WINDOW = 16155;
        301: PLM_AUDIO_SYNTHESIS_WINDOW = 14548;
        302: PLM_AUDIO_SYNTHESIS_WINDOW = 12980;
        303: PLM_AUDIO_SYNTHESIS_WINDOW = 11455;
        304: PLM_AUDIO_SYNTHESIS_WINDOW = 9975;
        305: PLM_AUDIO_SYNTHESIS_WINDOW = 8540;
        306: PLM_AUDIO_SYNTHESIS_WINDOW = 7154;
        307: PLM_AUDIO_SYNTHESIS_WINDOW = 5818;
        308: PLM_AUDIO_SYNTHESIS_WINDOW = 4533;
        309: PLM_AUDIO_SYNTHESIS_WINDOW = 3300;
        310: PLM_AUDIO_SYNTHESIS_WINDOW = 2122;
        311: PLM_AUDIO_SYNTHESIS_WINDOW = 998;
        312: PLM_AUDIO_SYNTHESIS_WINDOW = -70;
        313: PLM_AUDIO_SYNTHESIS_WINDOW = -1082;
        314: PLM_AUDIO_SYNTHESIS_WINDOW = -2037;
        315: PLM_AUDIO_SYNTHESIS_WINDOW = -2935;
        316: PLM_AUDIO_SYNTHESIS_WINDOW = -3776;
        317: PLM_AUDIO_SYNTHESIS_WINDOW = -4561;
        318: PLM_AUDIO_SYNTHESIS_WINDOW = -5288;
        319: PLM_AUDIO_SYNTHESIS_WINDOW = -5959;
        320: PLM_AUDIO_SYNTHESIS_WINDOW = 6574;
        321: PLM_AUDIO_SYNTHESIS_WINDOW = 7134;
        322: PLM_AUDIO_SYNTHESIS_WINDOW = 7640;
        323: PLM_AUDIO_SYNTHESIS_WINDOW = 8092;
        324: PLM_AUDIO_SYNTHESIS_WINDOW = 8492;
        325: PLM_AUDIO_SYNTHESIS_WINDOW = 8840;
        326: PLM_AUDIO_SYNTHESIS_WINDOW = 9139;
        327: PLM_AUDIO_SYNTHESIS_WINDOW = 9389;
        328: PLM_AUDIO_SYNTHESIS_WINDOW = 9592;
        329: PLM_AUDIO_SYNTHESIS_WINDOW = 9750;
        330: PLM_AUDIO_SYNTHESIS_WINDOW = 9863;
        331: PLM_AUDIO_SYNTHESIS_WINDOW = 9935;
        332: PLM_AUDIO_SYNTHESIS_WINDOW = 9966;
        333: PLM_AUDIO_SYNTHESIS_WINDOW = 9959;
        334: PLM_AUDIO_SYNTHESIS_WINDOW = 9916;
        335: PLM_AUDIO_SYNTHESIS_WINDOW = 9838;
        336: PLM_AUDIO_SYNTHESIS_WINDOW = 9727;
        337: PLM_AUDIO_SYNTHESIS_WINDOW = 9585;
        338: PLM_AUDIO_SYNTHESIS_WINDOW = 9416;
        339: PLM_AUDIO_SYNTHESIS_WINDOW = 9219;
        340: PLM_AUDIO_SYNTHESIS_WINDOW = 8998;
        341: PLM_AUDIO_SYNTHESIS_WINDOW = 8755;
        342: PLM_AUDIO_SYNTHESIS_WINDOW = 8491;
        343: PLM_AUDIO_SYNTHESIS_WINDOW = 8209;
        344: PLM_AUDIO_SYNTHESIS_WINDOW = 7910;
        345: PLM_AUDIO_SYNTHESIS_WINDOW = 7597;
        346: PLM_AUDIO_SYNTHESIS_WINDOW = 7271;
        347: PLM_AUDIO_SYNTHESIS_WINDOW = 6935;
        348: PLM_AUDIO_SYNTHESIS_WINDOW = 6589;
        349: PLM_AUDIO_SYNTHESIS_WINDOW = 6237;
        350: PLM_AUDIO_SYNTHESIS_WINDOW = 5879;
        351: PLM_AUDIO_SYNTHESIS_WINDOW = 5517;
        352: PLM_AUDIO_SYNTHESIS_WINDOW = 5153;
        353: PLM_AUDIO_SYNTHESIS_WINDOW = 4788;
        354: PLM_AUDIO_SYNTHESIS_WINDOW = 4425;
        355: PLM_AUDIO_SYNTHESIS_WINDOW = 4063;
        356: PLM_AUDIO_SYNTHESIS_WINDOW = 3705;
        357: PLM_AUDIO_SYNTHESIS_WINDOW = 3351;
        358: PLM_AUDIO_SYNTHESIS_WINDOW = 3004;
        359: PLM_AUDIO_SYNTHESIS_WINDOW = 2663;
        360: PLM_AUDIO_SYNTHESIS_WINDOW = 2330;
        361: PLM_AUDIO_SYNTHESIS_WINDOW = 2006;
        362: PLM_AUDIO_SYNTHESIS_WINDOW = 1692;
        363: PLM_AUDIO_SYNTHESIS_WINDOW = 1388;
        364: PLM_AUDIO_SYNTHESIS_WINDOW = 1095;
        365: PLM_AUDIO_SYNTHESIS_WINDOW = 814;
        366: PLM_AUDIO_SYNTHESIS_WINDOW = 545;
        367: PLM_AUDIO_SYNTHESIS_WINDOW = 288;
        368: PLM_AUDIO_SYNTHESIS_WINDOW = 45;
        369: PLM_AUDIO_SYNTHESIS_WINDOW = -185;
        370: PLM_AUDIO_SYNTHESIS_WINDOW = -402;
        371: PLM_AUDIO_SYNTHESIS_WINDOW = -605;
        372: PLM_AUDIO_SYNTHESIS_WINDOW = -794;
        373: PLM_AUDIO_SYNTHESIS_WINDOW = -970;
        374: PLM_AUDIO_SYNTHESIS_WINDOW = -1131;
        375: PLM_AUDIO_SYNTHESIS_WINDOW = -1280;
        376: PLM_AUDIO_SYNTHESIS_WINDOW = -1414;
        377: PLM_AUDIO_SYNTHESIS_WINDOW = -1535;
        378: PLM_AUDIO_SYNTHESIS_WINDOW = -1644;
        379: PLM_AUDIO_SYNTHESIS_WINDOW = -1739;
        380: PLM_AUDIO_SYNTHESIS_WINDOW = -1822;
        381: PLM_AUDIO_SYNTHESIS_WINDOW = -1893;
        382: PLM_AUDIO_SYNTHESIS_WINDOW = -1952;
        383: PLM_AUDIO_SYNTHESIS_WINDOW = -2000;
        384: PLM_AUDIO_SYNTHESIS_WINDOW = 2037;
        385: PLM_AUDIO_SYNTHESIS_WINDOW = 2063;
        386: PLM_AUDIO_SYNTHESIS_WINDOW = 2080;
        387: PLM_AUDIO_SYNTHESIS_WINDOW = 2087;
        388: PLM_AUDIO_SYNTHESIS_WINDOW = 2085;
        389: PLM_AUDIO_SYNTHESIS_WINDOW = 2075;
        390: PLM_AUDIO_SYNTHESIS_WINDOW = 2057;
        391: PLM_AUDIO_SYNTHESIS_WINDOW = 2032;
        392: PLM_AUDIO_SYNTHESIS_WINDOW = 2001;
        393: PLM_AUDIO_SYNTHESIS_WINDOW = 1962;
        394: PLM_AUDIO_SYNTHESIS_WINDOW = 1919;
        395: PLM_AUDIO_SYNTHESIS_WINDOW = 1870;
        396: PLM_AUDIO_SYNTHESIS_WINDOW = 1817;
        397: PLM_AUDIO_SYNTHESIS_WINDOW = 1759;
        398: PLM_AUDIO_SYNTHESIS_WINDOW = 1698;
        399: PLM_AUDIO_SYNTHESIS_WINDOW = 1634;
        400: PLM_AUDIO_SYNTHESIS_WINDOW = 1567;
        401: PLM_AUDIO_SYNTHESIS_WINDOW = 1498;
        402: PLM_AUDIO_SYNTHESIS_WINDOW = 1428;
        403: PLM_AUDIO_SYNTHESIS_WINDOW = 1356;
        404: PLM_AUDIO_SYNTHESIS_WINDOW = 1283;
        405: PLM_AUDIO_SYNTHESIS_WINDOW = 1210;
        406: PLM_AUDIO_SYNTHESIS_WINDOW = 1137;
        407: PLM_AUDIO_SYNTHESIS_WINDOW = 1064;
        408: PLM_AUDIO_SYNTHESIS_WINDOW = 991;
        409: PLM_AUDIO_SYNTHESIS_WINDOW = 919;
        410: PLM_AUDIO_SYNTHESIS_WINDOW = 848;
        411: PLM_AUDIO_SYNTHESIS_WINDOW = 779;
        412: PLM_AUDIO_SYNTHESIS_WINDOW = 711;
        413: PLM_AUDIO_SYNTHESIS_WINDOW = 645;
        414: PLM_AUDIO_SYNTHESIS_WINDOW = 581;
        415: PLM_AUDIO_SYNTHESIS_WINDOW = 519;
        416: PLM_AUDIO_SYNTHESIS_WINDOW = 459;
        417: PLM_AUDIO_SYNTHESIS_WINDOW = 401;
        418: PLM_AUDIO_SYNTHESIS_WINDOW = 347;
        419: PLM_AUDIO_SYNTHESIS_WINDOW = 294;
        420: PLM_AUDIO_SYNTHESIS_WINDOW = 244;
        421: PLM_AUDIO_SYNTHESIS_WINDOW = 197;
        422: PLM_AUDIO_SYNTHESIS_WINDOW = 153;
        423: PLM_AUDIO_SYNTHESIS_WINDOW = 111;
        424: PLM_AUDIO_SYNTHESIS_WINDOW = 72;
        425: PLM_AUDIO_SYNTHESIS_WINDOW = 36;
        426: PLM_AUDIO_SYNTHESIS_WINDOW = 2;
        427: PLM_AUDIO_SYNTHESIS_WINDOW = -29;
        428: PLM_AUDIO_SYNTHESIS_WINDOW = -57;
        429: PLM_AUDIO_SYNTHESIS_WINDOW = -83;
        430: PLM_AUDIO_SYNTHESIS_WINDOW = -106;
        431: PLM_AUDIO_SYNTHESIS_WINDOW = -127;
        432: PLM_AUDIO_SYNTHESIS_WINDOW = -146;
        433: PLM_AUDIO_SYNTHESIS_WINDOW = -163;
        434: PLM_AUDIO_SYNTHESIS_WINDOW = -177;
        435: PLM_AUDIO_SYNTHESIS_WINDOW = -189;
        436: PLM_AUDIO_SYNTHESIS_WINDOW = -200;
        437: PLM_AUDIO_SYNTHESIS_WINDOW = -208;
        438: PLM_AUDIO_SYNTHESIS_WINDOW = -215;
        439: PLM_AUDIO_SYNTHESIS_WINDOW = -221;
        440: PLM_AUDIO_SYNTHESIS_WINDOW = -224;
        441: PLM_AUDIO_SYNTHESIS_WINDOW = -227;
        442: PLM_AUDIO_SYNTHESIS_WINDOW = -228;
        443: PLM_AUDIO_SYNTHESIS_WINDOW = -228;
        444: PLM_AUDIO_SYNTHESIS_WINDOW = -227;
        445: PLM_AUDIO_SYNTHESIS_WINDOW = -225;
        446: PLM_AUDIO_SYNTHESIS_WINDOW = -222;
        447: PLM_AUDIO_SYNTHESIS_WINDOW = -218;
        448: PLM_AUDIO_SYNTHESIS_WINDOW = 213;
        449: PLM_AUDIO_SYNTHESIS_WINDOW = 208;
        450: PLM_AUDIO_SYNTHESIS_WINDOW = 202;
        451: PLM_AUDIO_SYNTHESIS_WINDOW = 196;
        452: PLM_AUDIO_SYNTHESIS_WINDOW = 190;
        453: PLM_AUDIO_SYNTHESIS_WINDOW = 183;
        454: PLM_AUDIO_SYNTHESIS_WINDOW = 176;
        455: PLM_AUDIO_SYNTHESIS_WINDOW = 169;
        456: PLM_AUDIO_SYNTHESIS_WINDOW = 161;
        457: PLM_AUDIO_SYNTHESIS_WINDOW = 154;
        458: PLM_AUDIO_SYNTHESIS_WINDOW = 147;
        459: PLM_AUDIO_SYNTHESIS_WINDOW = 139;
        460: PLM_AUDIO_SYNTHESIS_WINDOW = 132;
        461: PLM_AUDIO_SYNTHESIS_WINDOW = 125;
        462: PLM_AUDIO_SYNTHESIS_WINDOW = 117;
        463: PLM_AUDIO_SYNTHESIS_WINDOW = 111;
        464: PLM_AUDIO_SYNTHESIS_WINDOW = 104;
        465: PLM_AUDIO_SYNTHESIS_WINDOW = 97;
        466: PLM_AUDIO_SYNTHESIS_WINDOW = 91;
        467: PLM_AUDIO_SYNTHESIS_WINDOW = 85;
        468: PLM_AUDIO_SYNTHESIS_WINDOW = 79;
        469: PLM_AUDIO_SYNTHESIS_WINDOW = 73;
        470: PLM_AUDIO_SYNTHESIS_WINDOW = 68;
        471: PLM_AUDIO_SYNTHESIS_WINDOW = 63;
        472: PLM_AUDIO_SYNTHESIS_WINDOW = 58;
        473: PLM_AUDIO_SYNTHESIS_WINDOW = 53;
        474: PLM_AUDIO_SYNTHESIS_WINDOW = 49;
        475: PLM_AUDIO_SYNTHESIS_WINDOW = 45;
        476: PLM_AUDIO_SYNTHESIS_WINDOW = 41;
        477: PLM_AUDIO_SYNTHESIS_WINDOW = 38;
        478: PLM_AUDIO_SYNTHESIS_WINDOW = 35;
        479: PLM_AUDIO_SYNTHESIS_WINDOW = 31;
        480: PLM_AUDIO_SYNTHESIS_WINDOW = 29;
        481: PLM_AUDIO_SYNTHESIS_WINDOW = 26;
        482: PLM_AUDIO_SYNTHESIS_WINDOW = 24;
        483: PLM_AUDIO_SYNTHESIS_WINDOW = 21;
        484: PLM_AUDIO_SYNTHESIS_WINDOW = 19;
        485: PLM_AUDIO_SYNTHESIS_WINDOW = 17;
        486: PLM_AUDIO_SYNTHESIS_WINDOW = 16;
        487: PLM_AUDIO_SYNTHESIS_WINDOW = 14;
        488: PLM_AUDIO_SYNTHESIS_WINDOW = 13;
        489: PLM_AUDIO_SYNTHESIS_WINDOW = 11;
        490: PLM_AUDIO_SYNTHESIS_WINDOW = 10;
        491: PLM_AUDIO_SYNTHESIS_WINDOW = 9;
        492: PLM_AUDIO_SYNTHESIS_WINDOW = 8;
        493: PLM_AUDIO_SYNTHESIS_WINDOW = 7;
        494: PLM_AUDIO_SYNTHESIS_WINDOW = 7;
        495: PLM_AUDIO_SYNTHESIS_WINDOW = 6;
        496: PLM_AUDIO_SYNTHESIS_WINDOW = 5;
        497: PLM_AUDIO_SYNTHESIS_WINDOW = 5;
        498: PLM_AUDIO_SYNTHESIS_WINDOW = 4;
        499: PLM_AUDIO_SYNTHESIS_WINDOW = 4;
        500: PLM_AUDIO_SYNTHESIS_WINDOW = 3;
        501: PLM_AUDIO_SYNTHESIS_WINDOW = 3;
        502: PLM_AUDIO_SYNTHESIS_WINDOW = 2;
        503: PLM_AUDIO_SYNTHESIS_WINDOW = 2;
        504: PLM_AUDIO_SYNTHESIS_WINDOW = 2;
        505: PLM_AUDIO_SYNTHESIS_WINDOW = 2;
        506: PLM_AUDIO_SYNTHESIS_WINDOW = 1;
        507: PLM_AUDIO_SYNTHESIS_WINDOW = 1;
        508: PLM_AUDIO_SYNTHESIS_WINDOW = 1;
        509: PLM_AUDIO_SYNTHESIS_WINDOW = 1;
        510: PLM_AUDIO_SYNTHESIS_WINDOW = 1;
        511: PLM_AUDIO_SYNTHESIS_WINDOW = 1;
    endcase
endfunction
